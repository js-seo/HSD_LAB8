module my_pe #(parameter L_RAM_SIZE = 6)
(
    // clk/reset
    input aclk,
    input aresetn,
    // port A
    input [31:0] ain,
    // peram -> port B
    input [31:0] din,
    input [L_RAM_SIZE-1:0]  addr,
    input we,
    // integrated valid signal
    input valid,
    // computation result
    output dvalid,
    output [31:0] dout
);

  // peram: PE's local RAM -> Port B
  reg [31:0] bin;
  (* ram_style = "block" *) reg [31:0] peram [0:2**L_RAM_SIZE - 1];

  always @(posedge aclk)
    if (we)
      peram[addr] <= din;
    else
      bin <= peram[addr];

  reg[2:0] counter;

  always @(posedge aclk)
    if (valid)
        counter <= 6;
    else
        counter <= (counter > 0) ? counter - 1 : 0;

  reg[31:0] accum;
  always @(posedge aclk)
    if (!aresetn)
        accum <= 0;
    else if (counter == 4)
        accum <= dout;

  wire mac_en;
  assign mac_en = counter > 1;
  wire[39:0] cin = { accum, 8'b0 };
  assign dvalid = counter == 1;

  xbip_multadd_0 mac_ip (
    .clk(aclk),
    .sclr(!aresetn),
    .ce(mac_en),
    .a(ain[15:0]),
    .b(bin[15:0]),
    .c(cin),
    .subtract('b0),
    .p(dout)
  );
endmodule
