`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZM5xuMjGt1MYsF/EqGL7kiYV5dWbJJUBW4K1sdV4ct/Hjz60yl9SjjPLLOBo7z1JjlTYNB1eYrc1
mtItFpyTJw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J+1JIuunf3n83xj4btPG92Mrj4UkJWfESqPO+NKqWnsGbdF1QCHl93QiLE5wpjFDklIQlTxNWx8r
IigjjEUNH3zzb9/UU+CZa8forSmH3FZny6t8oGWpHw4XOiwE8QpaA1bCXx41UCdJviCY+KYTpQEB
1gnxRmAegARmYhnd0Lo=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
af96WGBLlfeYfBBoCyk18+mj7VnjX7uyGWyBMvdDo29BvUJ9OPtIOquP+hpOzT4wcD7SEOxMmuvh
vZQb+oNbqgusTage4+JqoOLi3oRpCXZhS+gBkaKWVCFj8EfccKZpnum/klvVrNOGl01VAY0wKz7V
sHCOV0agSbQNIcN+NTs=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k1jHUBokF0aLTHnZCQ+Ls1Y59IiYK+cq/6GoiobdhquF35TNOQIDZvs8PozVLLXigZpQfqgYT9gx
g3ZtR7zzx50IyyDVWQd+8Q9P1aVZVWjzqSkw0j5Z30NnDCZHHc9fGkj0MLzL1esdrbXneQ1s5mc7
O/m7ZTvPaaSXbReQMDlpRZWhcfIWDSzRYW7jrIk1rU7oTqxx+zdNjqLiRyQ8KtSE/Yq6GOj6MLaT
9hMu8L4/SvT0dW9gw19soT5TWgBiju7xnKoHsJEHFkrQp75jPuGxhAux+GUc4jL9wBVhT20rz/Kr
BMM78K76W5YTl7Q9FdcpJae6ydBm5WhWcW2+Pg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X7ivdX+Xa2Vxzx7eSFNgRwA2xKBMou8zzXf5TsaJ8m8HoReqLa1U55WBakDirw8TMs+RZebxF3rU
MDUCgUxoAjHUgDxruRmeCkWcGLt+aHBuNsWKhvhDefsNXlxJG8HLATmd44kd/dn+zGFpNTYB96QT
vXOCsRMA0+zCspCWPO6ojQgo+ubMf9AoUcfB5gxgH1/X2dd9VjxlAnav03ErIdjasXyL096Y+Ocj
C/p/Z03WG+T7v2QQljrmxBpfgfz6lzHRR2lph952rYU6JV4LEo6NJtQ0kP4596/CEAWotnD0Q6hh
3EHYhkHVRi+q1GoJueWVBaZw+hbKcegclCa8/g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F7v51tBmpmS3nIYzM3UiY61kS0qYs8ea092VJC2Rc/ZSS/DRru2lCGgqNaIhePgAScZ/JNFr5SOr
V/RF2ni3q86lyrQwa1XEmBnHgVAF2ap6C4F9w3Oxpr0cxhBoDNPq1fE8z1PjVD2qAjpbOPl7IdXB
z+9CRHq60XR1oPmbbjwerB4T/+bvFyY5SIHSh1bwPm65x4fUVhRnm5KOQZYXi6lWuvpI2QsKyjyR
jkoUx4X4lgzILXacFY5DJJkTShrHUmOyoDK0nv3PBka2rmrkMN/eYlrp5RojkIYXYBzettEfxwIN
Rt2ON5nUWAa+6YDUWO4FwnmsPZ7tre1E714HLA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 96624)
`protect data_block
G7cr3ww+abXM9j4X+/vygQmPN3LlkDCNzmduXyBzqJKeI4rY/VezFhCB2MFfAuDlgQnXTJqRbFdN
LToQExNDfQWCkxMZGbZxVmcX/1TwpPViSBogTAUh3zJq8MYorq5yve+LtRpuK4QeDVBNMm6qjix2
6B9ymhHJ50xZBYgTpOLcWPEiQI/GAyQIp8Y5tlVlgMu5P5t5qAJoIi0dtQ5M3r0thSf9AKqKiBTH
kC2YoCotJSV7uuCe8nqqNyD9kwQX2lbH6UemSYMiv18wldSZHLjn/CTATRqLLoIbsZGTcSt8OwL0
r+V5MgN/eVtFXNyvy1DBKiQVrlvahfcGpnMghjpfYn4DEqr3eJpVaAXNbDkIG/Fuaz2/YqyTkMeU
mjNtgFYsWL1GFM2J7M2M2EsV6DViqPj/lg2Z9rbeLGWpUrzi2cXWtTj+2srIRolQgpvoObThA3yW
cBICSFavJSHrSZtV/KbcMZhZx00SiAI97KkIL7W6MwNyePxoM4jFV2GuhzzfJMpMVrrOeyV6dJGc
NsJzf/ZTlWjEXNmuK7rqXjKbFIAvJlxFxmi6vtoaKu6Ms3nHHwkdiTGI6/liMTG/fSkiZ8QyQKI7
Plb1DcJaV3uw8ojm6KZd+ogLCV2rTuYxl+pJiem8lDOZtJqAjgkEiXx+pIxsCWLTQJ6oa9clcPKg
Yq5Xdtelt8xoGo3RqTZ6NnDltIr/SghmB9foNp2qZgjn/lhbPa7iHpWGNcnH/TKsKJ5ig9w3duwK
Sw5MiS+ggzbZu2BBDA1VewrUrmY51IelOK0WBwWctltSnPYdey4DFd3NBOfFvUQOm2bj8N4ZfTZy
ZKJGD/3moircLVnfHmKsfoYB9T0eYGa22u6BsDXNxtBF2OWxNpobwsK8dgm+RRVKqAKn7btPgnl7
aQSjJr6/e4OqHF5qRRjIQ6OEbO8idP1XntgQ8Lzy9obBEy3ENHvOd4eucuSFb30B9epnUzL8ZIU1
1iyTbLMfv5AGDwmCpL4mVYWjwiHZ9loJaKAWxIuxgo175rMq65feEsadtBNvrJV0P3Uq/2gwgzEI
OigkTKduIfTCtZuFofht1KyHERXPByIOF2OWlm4kXOfzPu0mrF1e/L2bsBPHFNlqnChw4c7x+peS
MAmFVCEfaVyOByOGmJcFjwLqAF4Kliv9MYQOT6QEyqa6crW67Qio55vxMS9o8EBee5Lm6jyAZQjc
SLU6CmVN0CEG0iePtXa3pi6rR8JBv6/9kyn+rKOzY/UKA6Gmfd5S3zN1iOwqPDQoF8y2Cq1QSJgO
2iyRpr1e3BES+upjXdyQXFM9T0xoL/ZXGMhpVYWzDTPonbao4xCoGwKlz/rztD0hp2BpgcDZOOri
jMZokPWzhkX7Abh+RF+7jbZn8C/bYi7/mZvbMm3qpIXVGyJufSlcD7eIffgSoR133Q9Xg1lK4b3M
0brHIZCRgHw/Iv9dRhLiPbFX/bIIWuPhRSwsOqbZAl/I0FR0XfL5JviXG8oqp2g/kxa73oUIKhkR
NXkANYDuzSp/57fmscsnSdlD4RfEBYd0x3hQ3tG1C9GX9a+7XLy/crBUuhbSqFEAnL3R7985yDjs
PdsCTr6JUs2CV/JsF4fAXrMziotlLR38vnvoI9B4erqglK/sI0grsQCscpLgGpOqx6ElmhJl1RyX
xycI5bDbBBZYKWiiWPeYIv8ApJ548PDB21xOeknYXFGo86HasVHHesxEJskNhZ1WrKjizW67/R8i
CxkdwB9XNjBWWVZJg2yi4mHRKz25WQO9jx9VLwYqGjLucflRSVGG5l+B308LsRrlW2D5/anv+O5A
sI4PAsvWMtdWsG2lllPHNLngNqMkRiKJtHQIoinJPbn1V8EEQO5pFNODK1POzMAfj7WBYy8KYEk+
j+9XYaX3lMym903IgQWGvSiXOfTAyvQjCIoy/l2flbeQgcvV+N+LkaL+bDd6qLjY3tFDToxLtp5t
23EHUVsSuuU+7vLH3wEmZ4HhhQ4+xF3l/hEmrOTsCob3IdB0wG02DavWVEa7PCy2Gt5AkuVMG0UD
w0tmZvZi5f1uHKZq5daYqW9xiFqgQaz6a7PPie9dJV0/7H4L0em5MTcmnkiOYZLl2KjEztRHtfOm
5BwJ4S3Sbi1Cn8mJnp1HF0Qd2GB46Yw6ZlErDI0cDLexXAXA6sxj9Tj9zXh3FE9/G5vUL9gWpMuL
zg41rzqYbyienDPZkRTXv8kHrQ0TqPf2vEcvd1vJmH63EqNw/8lRcgPjRUC3LTwWJ07RGl3a7PG2
KZezEJeKdtY2yZr6LUPv+aSF4TSMx5RN84/ZfWqmRIOZxn1rEtOzhYac4VbdwQ1wER9JID7wAtk8
qXh6N7RYvwkfqFyjsF2P6nfR6VqK/rtxZacpnd+qu1oKhHYYj66bcqu+Uaq1s/qsMt9xjQ2RkTMP
86SnEOHHlWJEOJRXe8hfICn/epYHrrmcQZ2T8c+mhEPEW0TDx2PmZKC2rI6mEN1iognkJvSV6lpS
h+NOtZV6e3AWjeHXCoRTzZnRnN329Ds5O10w7OVg0MJ2TUIp0UQa74LGTBW4bBEF6Zpfu+hFlgr7
dFYKrB9oHPlQtoCRh1hw9Ev3QNGTxAOJcIL37LPm3FuBXG6eeKXGoa106QFuhuicGFceZ8LkBTQi
tcZMHOUKDliyHAm3XM+91she3G8iivp/kGV8ittK6uQxRawvD9GFj7gIr63duC3N5Qql7PDh4jQR
C4B7Ga4FSlCrZkTHPAzr7yHEi11PHc4u2j3xcxR22B0m64gsSAPcH91G0fsJHx9oO4lRzp8ARhGm
xVFk6utgcpzITt2toTTBQODS8E4fgB6ERqE3/HiRM4GFBIS2L400FB+A1Tk5CCpOyaJYrBeCkHbV
i0Fo/EPxiIkQr5PqpKQ0UaJjn4fvwn0YJBvHq14slQc1+jauLe1FATDnphlsqh3+fHJYI6Bp5sN0
PFqt/bdd7jmSc3tcJ059j+kSoifaiYT5odUhf5vAk4xy/hmhAMt/ZHVAZ2d0o35OHk9z+tAt077h
RkSr+KJ58y3K6BugYO7iBsz0vlFjZ6x7V4ixXILPHU3vvJXqMceYhAuKYsI56+h+EvZd9Vxj0nKr
EDqjaF9jtJh+mbgF/+RTSrDAlWNM2LTnZItWJXYWHayYaqc9NPH/YEn3vin0vY+XZYnSRCpWUTor
Ak7XQDAkrzWGGUDeYsLFlUCAlDFSnE3I8laFMXWCOqbf7hzLOdwTEJ1Qm8fKCz3zbJ52ktU9cJHS
BMuGvE+jNT1FKxNpBnW3NyCDEaV7KjAcdfRSz1XCzEI9fgCg21au+wJPpREtzyBao0y7h5WxVUfX
5CS74TbEimdUetJWUSwtjuxrqAmroicjkC4Fqimc6JxUNuTRPeh/eczGT+61aR2XDPmAywE4Y7UA
TNp21PCAEMashc9280iDiV5F2ftKI5kpAJzubfawhadx4G99A1FziWkweQB+JI8laBfO67gHtfdS
rlhf/JIp4tlz49YyOJyFVAGtyHgscCyhNfHhZ+9mfcxaBvUFyuYaSibM3a6EZ6dk1ZfLjG6fOgGD
6ZeazMJI2MGpmDk4Q3WNcU+97YB6F5DE1Yw78BettEvLz7x2YNcC5eVyuS2HHDXUjuLvr+/jMMQo
oJUOww16NiC/HNnLxJdDc5DP9wdQMzFlJdGwWubLrK7yY6eYfjAEq5u4kjuZCv2ZDQVzf7wY7iaw
tPbVyKneTlvO5eDiXMbGTpkf03SsY6l6AjuMUlIQsj1sl0rMC4wR510iTSC7GwFj1v3LUUTP/Arq
v4+kkcipWDL20xfEGkE7fWLD+TP2zzXPzAij3w7vuxYAAiV0teRMblt7IkU7q/sedcjYNfBHOjC3
gFXEhz1Sn3/1VjQ7VwPaNymBXbNrzYg45Nh3HW1Ob62fo8me5bw0+mmdwcYfRCZCeFdQPoAof1H/
NQ0gMg+/M/zu3JPNIa38LfJhZ3mk/X+8yYDIRQUWWP4TIhqdGMt4cKl3FM7kZ3oivUwfNImv36t/
4AfJ3y3Bf4Y5ZHykLiQsWgdm/oRskduObmT3EOgHqmLFNMSSf3qfsgHry4zdvFJDezckzJ4ZW3Rc
5gw2JYIncl+5K/pNC6YaSU9W3kVSCCLBxdgFVU9PyYnLadux/GKwQALaNnbWgVnZrkOnaSr5KkoR
uhr2JeNS62n02Z/+pydXUdB39/q79Tne2hi2WZDK+mamvwHlS4GL3y47W7nyjVxwXtnjxupxF9BO
fPqZ26ESh/0hqp518FTv0WL2Wazwh40L3QMN6pp+FouDQw3ZPd1hyinGZBQNJ6D+IZNkQdkL8KrK
kxaL6S314quQ9CVuoMIAGF7jO7s1SdZdLKSXWf4T3tsaPhi6g0D2Ip80Gx5Fvkfd3fKo18IfFt2F
0hZvkiYfRtRx7MJFBC6I+Tldtnx7AsgRWIcRsYslMG0vnH1K+AM42ovF42orIWqMGcKzHPGZ13rB
NeVbG24IYsJJDt+TaWWWaPrPZor66hVf3KNCH478vIGk6/4Nsy19Cmb4FRHXlC24p0/+JF/myYqP
ztHsSf9L278Nt09ek00Q6smx1DcZSQ1KJM3uQljaw43yhs9WWvkk4gOE4cLObwblmAzGi5wxGvar
xQwSQGtBZZIuRK+qDhLTO3ql3bwEgLpWi93EKhibdhPuvTNmOtp0x3DsnuinL7Y+/M3QdLgVF9FD
0bKzFK2403M5T6quHC/rAEDEsd4URatQ8e+MIjeEh4iPl5SHOPhET2APpOwU8bDANstaH2KJbvE2
dG9GtZAYI08kc4BL1eOHVP8DGBVl5nyM75wd8K3riCP3Es1ChLFB5HKhyFvj3YzN/cQ3BV9LqtHj
SCcPeKWvARJhaqM2z3AzXOguNR7MOHnBjiKNrr3D/3GhFlJlwNBDXrAU+TXLtGX1H2noYzrhGcyC
XjJW/cWl08hF2foah+z5TB61L2LtESRr+DW+RclKorwaNUNzw+Ino5wgfM8LXDmvVUjB70yzCO99
QtRtuCASA+LHLZzAOBu4OHwM3cWiLq69tHLGh5wZ5V6R8C9T5fnNjn11oLzxaH43Ry4OvH75OJ11
Sl4Hkza2WASAKRaf9XN/iqGgb8dn8/M4riPZIK8AjvyyO6iwTJ9yTBbkjWHgs0R9EHELnl06rPIz
Ax63sUKtevMioxaFRa3eZP/337XlOox6+lGk3JMnXKhD5zEK92VxPN1CcMuB3ejaPBFk8zgQQMen
N+qbr94B53jgi74f3v3MCPDU4oYdTiH2GuakwiHoMatLkAa80UllkvITOmxWvRHnk1DEfJxoKGD4
WSPdCWHkfx5K40JNUkX7bL98muhpR5IVeH7HssCzuHeuUkVgAnljqOn/+Z5OQNeibcX5Gz6TJYQi
HHDAWORkSBPR4mgilfzeY0W7V7niPEvyiy6OabmeFM47Q0Ld9/X1LUUJ3baM4Ht7uwu2w0PQdJDw
OsMfp2fhrByH51E5jxvWuuYhyRq6xDS/CPkdrqgo4BQpSFYXUxCu+nVNDRCO9S8bsFCLeUQHBk7F
YBDRop1MGzlLcH2X8Ld0zIvWoGHnUBNj2kN/QozK6moElIS+QjFHdHlLvlF57peGFiyXL981J+9/
g+lcf5QspLYrvCkd98/adjy4bNbtql5gX4UalUTDnNi9sRUzj8p0WN/T2rMrRRAmZ5CvxwDgVjx2
H5vWGZFPhA3YfwZWP38yc2lkRV8Alt74zvGhq+jkyiwGUwrXCMro0rryy6fWJw7OV9s6AIDkT40T
sP5jD4oq3SlMLUtEgkt50OVKpHLpOjAXXeg+woV2kzTSkRoO8VuAZRhpnESYBYW1BiS3dSERl3JF
ZqOKmjVlf2DQiali4yh/jb3MFLzfRhw5zSFrpVaKAR6RO4HApWz0i/boKHDFV8ScwHy99iV/10bn
qx3+KjP/9J+tXp2U1Uk1ynpSCZuIJloCuIUWL1eqQXNgPPEubCeWtymGUs9dhxIXTTcePNpJjCWS
xKjzywPN6ywIFK8cRyFp/39dVkTCDaaYOWb5il9QhRtFuy6FZa9QRK9kGf6T+klF2cLxjAPTrlkc
l/CDHsENeCM+MnlYuvObyCH3iQ4T8X3fAR6HDiY0fMiJ0xh+KQPPuTqkoTdQ4e9j/JDE+s28bZA1
EVQAzAnlrUphAPVBBT9EGPDJha11E8UhQ1WDW1bwgNHiCMpE9ola5jGFzQYwmIU1ZZdP28IojPRG
cI2DSnEIZuyHIFzVYe6fFju3hfsebzV9JYgZbMt+witf83LFGnO3+ub9J3BaqU5PbqkwdXAX02Hy
2b4K4KaYVaFZ8TeFOlKHPLJFPq0RbH395USgITKvB5oE7WNRxnTHtjEJIHX5kWZoZc+pl4PVvOVp
pSK517Xo4igAdC9hfG+HE+d8rvxSKK4n+zkjd1F//3bxTM50OILBKPCphetI3Aq4qtTO94oDSYGm
OHu2sDr/Fns0LES2wQ+iADbeoccS1lrjHGiP/eDPxN39qRBA6JBJvo6+iniZogVvIr4VAAvucSJt
OF3hmvcLJOMN4hhrrW9iDv4Mimv+p+cSp3nBAjXew50LqdAus52SYF19lNW0JKx4tUbcn/QQHxUg
Rb5tAFy6P1BfRMYmjPPHZLcNAmoUlvDxorI7XHVXYoFv5lZvCT8kB6RBWyrNTdiuVgM7WBcfL4m+
jezlL+TR8R6x44msMpkPSVXcPnbKZIdf16N2kkoVoo0kK7oWl2GUUHvsyC+oCwvy9TjPjmy6E9zn
sx1N+qFI7QGydYVpKg83sSr6uEuTVeKbIxWKd8yIpIQeTPB7GibcrTYLaVo2qY1hyuYqr+SU2y4t
KIccuuSBHhnokTl6ljs584S0lj4ZFM+tHB+uZlt0tmVSbmHKWCkEQmfEwjyVKA9LDMUu1Odlsc7m
CiH13GGBZHph1XvT+FhKpYAMWPjIKI/3rz64De5NDEvrqVezAGCvd3pMhOArvLgGK4RNoFSjtB0L
QEasLs+G1VnXrHzzoaNHmlsZSp7qt55Hg7crEVURKtNloTIP9a9CCVvCDr4NZJ418arxDzXB441R
/f8CvE27E19SQjlhEnBpmbIKmzvnIRgBWVum5x2GZdHuK2brTxtjqBcWa142Rk2DtLX1eXwJE7ji
ZVfDkWHQpX2gweRIDe5FO9RDnuDI05XJkgkHio5zsjnLEYIVaxnra64Wyg28tOm6UmMfwWeFpyv8
gE4scXqHm25uuhx0Fv1YiMEcQ/BHXl6oa0C6aDDl1lguIlAuxmLZLAZgyWQAoyFjWNHHCHzUvA84
3JLgeHVpGJeH5XLXP6vR/wCWSGsXAQgBtCaDdxD/ulVght1a+9YagDBArt1CyjmSaSIRJA+RlyeO
+qE5VlU7RqCgnSXEQDfJcDmCdInQhDtyvZuAgwIla4JwgYqtz/ZIaBgh6ngjrKYOjtQtyeM8sq8y
L8wWY3sypLh+N3o/+niyBLNT3Q+fMVS+2CxPZt1at9QxouI+UMwPTyRugclrLlVQmzI0+0+8u1Jm
nIduXeO2HYN2EYihPiPlSLULRupvgpy2kZp8hSuiTzrQTbwv+aPA45rZihR/qIq7lOEK/JjcMiqm
++pUoOBvzG4XYhB0W6JUfMteUPXpbP+ly7mNAZEWTSbF5W5MtZ4st2/4r2WxCuZvWz6KXZwu5dZR
GPwUfN3Yd4CsyrIAscOJKqdQk81Vc1Hwxd9usfGv1QsCnv01KxR/Utx75KtNOSaY/QyS6lP1zfEW
XvhcvqCcWvAXDk6WZ0owSPFkyewVsDmSbesZ9NBOR/h/Jp7Y2RwIcBa7S1XjjXiDFBpDMo+CBL31
mY28tEO19NwDKFhV41AVusxtqtSFcUGORuxY0CbM8vQkeK8hPajPRksOyoXGiD2u6WCCwrm1c95k
m0Vna1eZCmOCt8vZlfBAcGI5rGzdv+fH5n8tpqATS/+bnoYlFgVekeQaa/OWD80ayMOZpNZdxWFH
jCdSwiFAyOqzUo9P2gGJqOslZaE3dnRdNiTa5d0NVssZa+/zUV0Gmls64DZ3YZGaLPQgeQcUQyuO
Ru85bSqi3x90RZ4IeAcVKKWcrFoQ33sgIYmWTcy/UE1x9BrDoGgk2vzzsPx5E591hs7QJChuW8lO
mUmhSw8aZ+S5TapzrHKgkj53PfXFNlpK3aU6PFbgbmqAtf3zR+aBQhjjKH5CG4dxeFE0XiTjg2a0
kvziqmXVFyuAZemHBWQzWuyxN9iNSelw0mQC6IuIYHd37aa+nMXaSl8nxlSCO52vaA+r2uSn8Gn+
lydzDUbX2r88PMRI86T7RyG7RD5ibm75yk/YAsQoLQENQg6QjEAcJlJOGTH4LB7BSTl/NlRXDeip
BuZ/OAnpXE6ynCA9ESO497y4xdZwgLvQdlc8Xm46LpzMlAnmPYcMxeMcM4h8kbEZumtDj/0cJBy0
j0WYzs7T7HL6yQos1igvJPkEOpbx2gfj9tlBG5H2yUcrZ6IEcHlMTUDom/d1uzJAGAiKZc77PN2k
doL/vQLdSDxm4QyXkSX6JeXfPHw+sU6H9zEU+rPGw28aexqn+MxOgXflpD9TP5VidvtyioZs1AW0
7wnnSPMZsOp14pv6pzj3E0xzyS99PkhvdI0J8mSOjBQgNFuqbdIlsVXGDgSJ80CtBXVoWWCrvkio
mZnsf8vua85qu0on0IGNozsvY4sbPWdgfJqRHY9f9+zhLJskNe6U704Pv7wL6TJrNSqUmh2i4JWs
EiT5A++Z8Do45P1oC5OND7YEPg48tUQw7FpvNepGVcvkjx8LJG7FKAFe56oFJsgTFpcZNxCN9GPM
2k/t4p3KtKF4CnWpfXrbo/2D0wvXLbwksMSaOCrum4qHxmhjIeqfT4+w523Jk4+ZyEvX2rPO1SbT
T6dUTLZLgXPjhqYkwAYzUqHq8IQGYDXOzIaWZqsTnvDI8wjArgbKBgG918DdiuWtjZdpePaDtdum
Z82ELw5MxGF88tvZ8JRnMSN/XVsdutJSPT3P+QpNPGJ/IlMzFngr3nADE3CsSBbtKR2VaWnEjLV+
8cJ2oYAPcdftF4vmwrYS9w3tz+tYBXLQTK5TpGclxKy33llygR8YgkWUkP7vz50vCG9owpj5Gb98
pedZa3U0KMw4gXV4Qvh1OGKHL//Kz5VMvmhyqMxrOIPiuVyO3peOE0TFoY9Ti9Y3Acx0cvb0MJvs
RJthiRX2BZhQGEdfC0xrUVodwCKIlby/zzqMUXQsKipRWw9EqJT2E3ENKyx7LyMyAJ/CsheQVge9
hH6Y8StiELGawWZun//SpUELrfSBgJ9JoO52EH0N/Oc8OdCBYzd9rq4JUq3M47zpA42OD5LOv889
W7092CtDnwereOn4KhrHiCUcYaGReMTgo6OopvgQzGaFj3DOpD4yGLgbSGIdrmwqUPSxjNbl5dSw
MDOyvEAMkASE69YGKlkqf+lv4Y3SFUx9ba9QkusFK/dh0t05iVMYhldHrT+6bBsHG3BAf9AFaqoA
TvzM4aZX9kl+7RPPKTgeTS2JplyJSqjR3tVFmmVcz0Em9juKn5y7tWWdb3obulw29Sh9QGPFtEGk
k+8JxmCmCKd32VxrGY6h8jWaSBh7bnid0KOT3tv7f5TFVxtsGG6mX5BCcsPd/Js4mO9pf7PIsxbG
Ziu3BsVTbZB3rh9OrIfg8AhBkJd97OszlA8YI7Z7xB3bMckdfuW6RWiUI/CAxmFhm9O/dUL4tzWZ
+JiISR74gmk2bG0Po03SZ9hI+VPeLT3DgL8H39vbFHl/ZWaS2mAt9LR8JoTaSheZWNSy/Fyxjg/r
9BZmHuunY74cn766ecqon5IFC2L4igIqPfQ6tpOS1ymC4zsLgFtSuO5eLy3YoS+PrkS/Qa/mq9QI
iwplXef0wqGgMjUhpnOZNtHdxCY+z8VliMWCxJBCPeZooaH4jvGvAfcWjWceR0tiUME8RkW2lbD1
BODgvaNo9zmGgMFYms4qXx4mH2eUoYKRi33H2ur1ATeducgiIUYNuBegl2/dt0yunH9BoUS8MH57
2gDSNEjWamaYCopZIKyBgKY8BIZDfXKq3Rg95/C6/bdl7+DC91CK7v6gDrfsw0EvIyWQv6CmZsat
XvahWiEHry/0IfUz/BzSCi7CjnHrw1XsaSJsd1keXDdgOkTY+G/OnRB3vVFIAJ6MvK9yaAB1ZZ4Q
wNPVhnodgM4x/uVxCYVTywEYX1Upp+UY8F+2DAraAYgSqsStuG5hMwOysa0eK+ZtbrUU+gE0fUTi
O4LOHtFgs4uYHFTlHP7VrgzAyYvPU4kor1WBS+gH+vg6fKIUSU+JZw7BozvBftPZmf3W7X2btH2o
TYFckbKASrj04Ltw2C2VDGMzgSRdlTQ4nnqJRp+qTYzQG0YCq0Nr6J1n55o0uFEmkXiY94DDBTEG
eB1Qe7kFqZtt59m9uM+h+oQKx8W9y5z8cy7LvcjXHHuf9S2UcZvW8auLjxzKahPIre0W4KQ4QQwt
BU0Uv9t79q1GTKQaM3LzXjNMwiL60lQT6fKGWDtR/EokWjcdlCIhJlYodN1vg6CTOcJRPSUJWPA4
0MLL6KERc995ifO2Imsg0PVe4clSAVDABdWHlTqKZKc0nsy6ssqlZ7G6/iJd/684b5k+/CFeu1dh
zD2MRuPoj6Yi4GScUqLOjwb16K5AS5g/Fx3b50kdB0qHK/7XKIayt+MakQ/I6TsBV5hkXNgcdXiW
gAASo+gQBDyoRReUDuKUZEOfUaAC/ASLzn1Y/Wx3owCxvZSpqWxrkjbCWo039/r4c+P7MLGdktlK
HB3wOJ0btTDJM5ncGovO1Cy9eVhH2uLy/viZYHusU/XP+FYWIvvWF1SR4sDvUdSUBStZl6Ku34rB
Vzn1Uk4jM5Y0evhF4UeqODawkbs0xd6xwqM/ISXeZOjUsPbKPVck/F3R3WMspBG+9gmMo9A+J9+j
3wkDvzKVejeKGWvO8jM22IQ6/I76DJkbGAOXtgDO2KZxp/wXvHpEAYAtO8O+N87RQPGCHfLklGp1
i4oPjdnsNCJuvuyOV0/0HdLCb1HcxIz1zsZXdw4dARZ2wm8KSLjzEmuWFmgBy3jQeCDQVvjbo7iQ
0KPxy3dBq0yghTpmlfVnASQy/FsZrL4CdvLxNaoMTLyaT3qzzIcejnd4tRFotXCCyb56yYXsicJQ
W1zqyEoioCy6zB5Sdmysq0+cFrVuD6+C4verytUk5PFOsr0qb3ZqpxQWSBedDDkU9YISL8riEZBQ
rN9jUF1XuvVDJHc4lUMidV/WPNKJJTijKhb9Zc73wcCIcrlhp9bvvMjWBuUGUL6+5sX45VQVaqvK
OHAtROheOh7hkqZ62M8JjcyB81sfFNZzvlhgHY/tWHPsXArm7MJr56qXLMYR5kHN5XVHWQYVxIhe
42+yNPcPqJ5OQD17H/oRgenS4obubtaAOR4XJA3t++sGimCumR95jlSoTvYimt5TYsgmJqcAnbqr
LT7TXfv8Ko6eUr/jTHNqAiDhToMyc845mLosX+I3+pnz8iGAC8qyJWSbn1+Kh2n7bdVAOYTR/jn9
v6BTsFzfvvMLCWLQNusuUeo4OMCr9CKcrwfEZhzZCNu5a+ZlFjlOIeru+VuBBrPWpOQxcE3gAWiE
rR+ByYQr8gnnyXipZhsYoEgAublM2aJOXTZt9IiFebSlSw7c9ReAafj5bjXwnYH8ueRFDSIrfWLs
cA3GBBbgNvA0cc5jE6kmU05IC/PQmxxW6zaCwSU11dWxc5N6hp4ocnLSOtKLHCMeH96a8MKAkxXo
/XkDJ7l2DjZheSjH5uQBPoWNr2teDRigZpcX8ZGEInvzOKV0mNnGe2jSFT54t6LSnUGJM4wobRcf
Tim0Ow5/+GQZQSONQASCNiK58ox8JEtlQOIJ8cUnAEuBeIZm41DJNi0699N5bDo7q8czS2UqZ5Os
g5Z7PupSAWaXlyYMv07ZeLQgWtmLnbzEAzv0yi/ipDa7B7MLAl95/oyRxstFZ5gQdcKwl+uxCNvz
m84wq2/A44l20sZR3NuXcoolx0HXctm/SlJrZplGnfkseA6EkdpAlvhDVT7K60cRaTGBQJdc6bm4
LehOOKo4G1PAkckL4MfQ0gjZyNNzf2hNbZ3qJojO/X95DnRfaeLuEcrTYGCfvzK6CuaVE3UK60Gl
GM7IvIirEeDzvd3w6ChME6YHiSshAmn0+2fvdjzUixAe7PHabOlJImpDM5RRzsqFsZFJvGUnKR0c
x3kn8ep6BvwYs/JNDkgn3ARzzJXDWUUlnffC4k/hyrVtwukgFcBPuu16rGo0Vm1sp9dfFJFdwesC
BhKXvDMrEpT2+ZX+Fx23NTavfZ36h/1EV8wNxlvcKztt2UuKwhfir+3EgJa8SdkexL2jYmxEjDoC
NQnggKlaSjFw6/Z/N6a/+0fA3ioIckgwj5Zhes0pualV+h00a1LRnn0AUrhQiIB4jh9uFnKMEO9F
5NpwtZEXoiQuGELm5fE9jf4j2QteynHjm9ZidfGNOyuDR18/AQlsA/BIZUukm+nQs/VUUnEK06Al
PyBjZTrmgK9PNQhQaC9bNjccdvJ0DhoGz3xbpzyYkApMVUFOQ/NlLmTrKfur7VnBN9c6mbJ4g9jz
Xr8JIrCZuNfcS/Bs4EAjYb83iNEf+0MU1NAk6xrLO8p/KA5SCNuGGZLzvF33itjjrlvR8P1Mcngd
28XUaUMuCIXjCHWNI8id+vaiSTj/Oa13qcPM/S1FbsM9Pwlt/nvtvCpN/FclkJJcrT6tfFK2VDc5
8OFk5dxDzNwjQCi7ceZs80EELVAyGpXTj5KJ1Fp48alQwcP9v00KY9OjFthokpdgIRSRLCLiW0/N
v2XK4nGCysnO6y/hSNERKEk1byT40yux5R5WZIVZnGDiKmTnWUAuHDJVBV8zhfcqZHJU143bxv0Y
GTVMfX/aOS0xx/qZ/612WSJsveRcrKyY7fRSw22+NQzhBlMDrXmNHC0WmWw26k2CUPlcxYsTgxx/
DJVd1bm33nHRme016AD6sYHtiEs2fy+T+ct6tLACEg0DCnhlH2PwR1/0pa7nysLVjzHpiU5kBJId
X+Tlgvptil8gbqIGc06NqKaPFzzoyT2lQcKXvSfIBjSplOI74Vh/iTsuZhtIngMVRYt7pNqNMSX1
lTiY0iD7WdzlChijyf1rPHvkagdvVoIMbgG6A4CwCfRO9Qr4KUL7iWC22NeIdLEVh8Qf5xYRJAWJ
qUY4osAC0IuHsaHdi/lm/7pP2JMtczUWRGV1D8l1nO+8Ws368Phoqg/swglex/UyJApmkp8JWisS
hIglRYwk9XRMswvlQNRzFMJXg6PfkpJ/JeMTb832aPq8cE+46/NvOLgjX3q62a34enBFNF+dSPGz
9WT/ucSTxEA96zyHMLw3bWMmhBiNnTdtmhZ3NALLMfRB3pLGPK+yNUGG6ZcLkk1+9YjKhHe0kTj7
cI10Yj+oihSwj/BGIRTHInTcFEI+zasczeshzWphRp2rH5il/Fn8vj2rue1SuUn+WAyDa+JZPYWy
XepqWrJNfSxLh+SRjS/OrRl+jQh/JJgHYJeUaKMpUVO7lDVEuZr8b6TodKpYp2GUNILT583+YDmS
58/U4NlVQLzWOnnXbVsOXGjY/svvRqSKTQOpCIGwU0wPm16JtDqfQZ0hHIwpdqkX0HShhIf4uBOa
HoBZtXevhCEPCZp4XOv6n02d0WaVi1wKY9BTGYxjQ/CchlNY3EcW+CGlIYNEWZ3ZgbFJKskVFnF3
40v54IBN9Ngy+muV9FuDOjmwHbhEjj/BPQRjkH07CSUT0Et0V8Wod03iPdjFqcW0JRZUAh0lv22J
mejSVdfpW7wdb7hM4ZVZh0n51UzOBVJ1GB2MTNg3XD2ZI9ZlwIXP6lH10qkYQ/Ic/bUqQRi9d3kj
TNZyvtZSmHDXGz2ph8E2SjPHh3T9cTHnKJ+AtCjUXretWUzwXpgho92ORIjd2YY0MIdew4bfCP7p
OLVuwgh3esr3sSwJLWZJ07QEhPkXV6HuLAOIJncaqgPRg2mM3Qd6XfjyPWxatQHYZcGFq7exLy9F
jdsi1E2GZ9EwncazaInbrDEU2/ykoAS/ImGDUm+Wsx7Ma6Twa87OLGJrhnqCGI/fguH2wDfyl48i
bsiRr3YfGrRPoCacYx21JI4jF/AQV48SHT0OiriOb51Qla6NzKUfnsrVldq4DEZAbvych2PcrlYB
tEQHhEmU4oBXjkVgy1I6GzfusxiIfk6X7VZU2RL2jHygvZslNwdBsQp0gFRAwaFSVps578gXeVkA
Ql1atIQLtNpRWdcc+i0apD0vv9GHkuh3FrgWExN5UYDOLCnw4+E/rmrLTpizEUtYRVCXC/HMA3IY
7SCQgsMRFsI/TZkWSe/GgLk2kn2C2MG/Q8A6br7RCQaxddVkkQIE47P/bjCT+GuVMUJ7eS5WfDkE
8Y/JcKcbYmgzk72ufyWOqpaHNop4tE+jC6Agqdyi2gr+jCTqM6c3nr8CwRWUJudoKL28BiJBijIK
mN1NBIBkb2C/zkMPSytr75vURmHRppHPFpJkPNIoA1qJINB55SEIgafrabQER29jUIHTceNZNAuJ
u6J4oxbE39EbcH/U2fWd+3YCNxMGURtJlTBO6J7FsngRsi+lhPa1yHI5uFcybs+wX0+Orpa38w/O
AuhXfGK8uX5doZ/U5GDK9GdxKUma1S938+2vmJ/dzkrQh8EnUb8Pw5JlxeL1oAd9b4SvI75FlRj9
jfYgsfzloTT6gAnbAhpayENdpltfDdgcssQ1PNDHbl+RxvV9mzgbXYntn6OIqWLRg2hfek4AWOj+
TVcvUnKXL/RE8KAp9cykz385hJTfsz6jWoEmZArBjcvSQfW1gmEByFsIaiPH+P9HY4P0IWWKqqDA
Fib7SelAnTFkoJTdBozB6b/w3XsHyz8jfQ7WIKKNTronIOSV1bc2gjrlwVD+deoSeLUGyDYg55P7
z+l5NidFb0K16Vk0b7z/kLpMAbap0gxUNuxftikJoGkOOEPFrXUwwZgN6vnXgU1bn/vOsVGh4SZC
CecqsGNILa3ouADIAqvAdBKb4aBsxwaoPwnqh5+3HWLSUld/17Zh495t+YFDqK92X4achftKnXiD
N4mh2vT+QK/tnvrWSOhBA2vF0yWUhUE5jqSH9tnuPqP7snTlqKUgDvBD2lmIXVmwjNJFHIyVsI7H
dZDhS1xxVYoj4UF+t0y2kvnDyglGL6g+ONJqj1KzAleSWhIRfMLuOcTKFvkf0PjCYY2HP5+DWtr/
VmsKbwdSj/ETLDq8fnE1Ts8x68sN9GlO7+VEYGtW06P49oYx0/7SRFKBRT3GjyMIJRCQMl1G7evG
CxBewYBTEWJUuePh2owdlY7af90kj1ow87uWNiJZxGO9J3MxDJoOdwnEkumrvpgM3uZ4IhDv96L6
8IeeoqdhSDiLPR8tyLukrGRrGVuGV8FniUEKaJk8s4/YZ5FeCf6cS47vj5ZVse0vDYF2SNthv9uL
3keeoUv8v7DWq4SRmAhzoRqiUMet+hCZ4vDx/JmndtexcKP24EmB+iLRbBywujTU2swB9sqspr3j
n+uPZEDJFqB6bW80W38LMdQFSeBjU6ry6zH9dNK3GuuzdM94VZmECQS1CZhzFq9wLEQG57IMNBKa
Q4lKJVBT5kPo9lKHNo2Sio/6zBUdLRu+ra3pe6ATmYM5YtiyLgLqMffSDw84gQ1laPWNmPmA080t
tjdftPZfNW5l7D71c5J0Za+Xh3TX+97EPRPyNnq/G4tBk8SnPaOXMkb5i7AlokplF5Dt65BHeDip
W3sLP/lBLiMCXmUVnHY5JUjNMoRhiyafKAP/34pBIr65+AkwEXUCYdmP9pwIDTjL+Pt0KxLM60Vy
6bUza3cLBjfmJTmvaRfKUuzn05viXDpDENGZVpBxanIoYzTYauVhwZsIUoZC4cV4Mxd8G+Glw/Pm
SRyljyPOeD89zzrEtB20TJeGsctb7zr9z8H1eyRByFxO6QHcfOs7aN96wzuK5saulgKZhj6ivk/o
Q4l21OotxHEwXOCXmDIMRb8j8m4NHGvmOmZihSW6indTnFVg3/nckfUnlLKlKJfATtqENwU5KQ+j
Jd1JjRUTAyLA5nuFHWUzmZb2CRN8ZY0ofDNEphqdvZu7coGO/TWedc0BUEmX9yaWc149GqCZ3Lb3
yePzAHh+ysLhFKdMB6XEH5XXOsDb0Oetvt+fbK6R6qXWgM+0oOlpRUJ57ePcfISnYb0xA7KrXhX+
pT8nW5tzsROwK9DHfvJCKwvEEufH3++shBK4Gi3uhREMDLOCwYH3DUjCZQtgYulneDpdht+gN16j
RaPxMsLKYnR9vXYr8AEd2t5A0uv7vRCgMuIEIvcjWjKutWgO/dfIDsWo0QpAcYsHNsEjoASPxf/a
XT/QfLcR2/2WEYO5Q9RfV4sfqGRNdeTPaKW1DAQQNYdEFXTWUH4tht8MsM5M5UKpOSeInUU2ly0h
mGYRQeCj4Qg1ht7o5oc6qIm6sIeFFfP7tXJweQ7Fp6m85l6HKIAr1oSDzCUqqGjCg+mgm/t2AE2e
O4NJAqiBm0tA2PEFcwpzZ3sBq5musZ631nEhbpcz+jPYT9tLLRyQA77rvh6bLerGJN1OuX6F3lZ+
LFIHRwM/C4w/3Y8ce1eF9WH8yQmq+mur+ZbSSwJeLiZW1k0EnSQyi33Js/Ely1e7pRWpoDCwmxXk
e0IYde3SGqVNJNXgKRIaJU5RMK2O8Fb4YmvCjG6nNh6EegDY3VRh/ngo3aK1eSJIDOfULoSaVulj
7vpPpv+YVY0LMuLDdIls60CDc83OL5Uoo/GnQw+oXsXvZKw+itP/zfTyCjzberF+7NxaTCCIT5AZ
yqRDEpDmpFkGnywjsLkoRJkaCFEHy8q7SzdYX+I0E+JWw9JK9EkGWv8eX0DuqcEWX/MCTUwHj0XJ
VaeXJ3cnJqVRrRRWV9HqTwayOGB+qV0JBd7yVbk8w0sDD2vXScVGCEaZgAErP8XVHx8Wdb2Tic+O
zXWWF8W61M5CyVb14b/lQlOxQW+YL3nDp9WNgMUe42GTFz01jJ6bYESqQv6fdd5/FsLgjeSCylIk
DK3AXE7bpQc1ODI8O5Bo1c9R+EHpAQ+d9Q8MEo/Iqp4dv2XDIdE3xae5I/xvpAEHdHZPs/sjfDc6
e5Z4qhvpCYtEqTDY/9q52G0E452ZX472DA/oww2VutdPvXtpQPfFQpy3dDcBQ1wZHFu1GI6YxiAl
ZeFk+xnH4+WtciQLVK9y9gvkEFX/jWwHLsmEFDdAJ+U6LZ6nxGOWndHU0R9X+zdgEDYF8pCp4PaV
P2e4VIlWGNKGBon7M1EYcAh6vT8ZDKT8rc9u8FM1pgIAJE1HkAxfYA+6addad2xA2TKUELSFXW+z
McrsSzndJp/CTgWhr8WvzLQuOZFu9FwwwawoIdKMYT6j+tZmxgwXpz9BHhP46mO9rszQ5nN6p+tR
0/mW2nXBgJpl6D8AmlGa5Gyh+Ojk+G1nXRW6K6TLc+Nt3SoYlMqgnvcnt4aqdd7JxB/fqcEuaYBd
RoAF2CMqLkGfvLhhOHSVhQaxT2xqp3cE1sOsnggi8NDn1PWQJmFWOg2SKoSyoE16qU+P/LAjWRDn
RNAIS5aXyZx9wrjLGwnUPAi4tjm4BMxqcq/051CTNPrsP+YNiT3fx4Z5JZJbPq44d4DkMslyyt0z
T+aYLAiwFNC/YzVbhkyFpUpeaAJv/Idl+Sot6cpO7b67+TilcVaWMVhK0QTLBMdSr3CnGh65pUNr
KRrLtWl0CbQkrBJRJwGXZycQhynvog802t4Ui8vhooEZ3Ex5e/BW8uCRJN6o65+/4KOF4lWFLPxp
CWyPOG7gNLkMF5bUbTw88mrK8C2A+km7Qp6szryCmRoXOhcshOEuuuR9BGqF/qFIyH0/IVPwQAVq
y0sRsF9ZGJ5nWLPDl58xTKHsSNYEc/jnkMxHEnaYkuswn9UN3AKsOmqhNXIM+sI7pEN1n1MBoQMT
5F3UYQTk9W0VF+cHjyJvlcoRNCgZBRpFvz0jw7ZwHTXiAfwP2ePSCzhKuK2WlBLZAP2TNdbG9nxD
FNvQJfxVfaLMhEkmLOaczk8QJekdw3zGZJdzFqTIE95rFWH+hu/CdG99/XK267A/xYFJ/2odqU64
ne4MxDR/y/UCL8NvXOuFkzpoCsGG5Z/DWu4qLwi+ugTK2EqsvYMmmyTpGBB+QLwjxEXhj5I8T3Vu
djEVxjtmFWYSghBhgnoVKwrthCDgdQNY7kNSLCOWm/aB+1sHzFj93XhB1d/JH5wKNTYbwQqzTV1U
iFEI9QzS/eE/jWfbu3JRG5TgiPGJj55ZBZ7LU8t6FiyyyrAXNIMBdanWPAtc2+/hE7483wQ+7lbz
/K+P4+Hw7OtBej8MtSvTR143ieO8KIjlZMLZlDo1oQA+ZzeEE9gGaQh/dIAXCW8+Gn686QIdUQ79
+q4Q7fJ2Gd6TxwRTM9e3ntmMK++8UYFaaJp7fEcn1TCVPkm79XR9wuMg1bXElJ9oCrxBl/YKYOPG
matQPJm/VDp9uprUsBWWD7HXJwZ8lyvxNH5rmv6GyRQ1iHuURCfg3tzOWyIHZmWoy34AL+HRzg0k
ZDSgqUn9Uqi/ZLdMmnKBVHau5A6YgFJXcOsg0vW7LLHGg33KRrGgzdJ+GfG2AdzIAIfCf1sRzV93
ghsgkZAgYpo5XmhiUe/LHKjpysSRY1OQZHDyLuPxVgS0Lk5OYCMfj9zzDizlIMqGeJk7eO/h/QAP
9R+rvg+wJSIXtt19aiT84RxiDX3chS9I1LnZo7b4qY3G6CR2yz3A8JmPHqELBE1EaW64B/o+mrci
hcq4nDSnBj7trKK+rHpOz4sxRrzz2VUjwnOV3hHM4ukIh42DNH0bBm5o+Xkq97+y1WJxgeEG5mOA
iwFnarOIRy6m9evyoYHKl4KHDq+EeEgDL4OesI41XNwHnM82zMMH3HF6f6CZ/uyl83Zsf97D/nex
S10NEu6CTpnbr/C63dZl/Tr2B+kKAfcZrCjMBIiK4hk5raJSimHlpnzmtSSEfeYrOOmilSiLaUDM
ZvhgVqx565moZEqG9mU8CMGhUk3VygQn8UyMex9otV4kJ9HwbKPkhBq5MRFKykeMAgiC7TxH6PYy
hmDGy0pGlcwjdq7R35nRg/RN6DrOKay88EIDKDuaNkc1dH6IV2ryBl2tdGXKlNgp8FUKuKZ0s+SM
6Er2PDOsgTf9+6+6cCnwjZzPctynWJvMbqhAL5hWt7aSN3oqMCoSlcfG39vsSoUj4NjEQn+cmJ4D
778DIeJ7mKKi2/E1Mx5yh3AzMJvK6tZwiI9MPF13NCODFXM/rLXaZUdiSaWQOu/weAvooMeZ6BiN
DkBTCPfiJ5lzvH2Gs/gNc0UxENCs9j4VKPR/WC38rDGmYUyvNTlmqQ892QE6yQbu6I9cewj63PiT
iRiMEvgCPvCKv4g97t2pXR1R3WfFEIcVO4JuTLBFtkRa9c3tCfR86iGTeVXACfMeqZRYOrq/0U/z
CGt0XLFNlLlnJkdv4ikqLQmSzUL+roK/zgcL3638XM1aVzflr/M7izKOAs90BowhPLCCHXlTfvv6
rXZRKMPWIYN1ba8XjygTzXZBkTLXixkrXnGevaMOnfBwmr/x5tID4ejz6JMynwEtbLzF1ZvddLVe
ix+BYuf/W0D5dIlryBZTQtxiVyrYDTnG/CoSEr5NMnGfy1SVQMgUeGx4ycnt+iATxd2MuNhF6+kz
WRnf6VYu0LhpQWQXVyVTO+1PZti+yg9N2iRAqcMaS8P4BU/h8NDSUnRwcEYimoS+L/DsJ8dNN8FH
Gxk9eeaT6K96xNUT92aIw4Gllxa1Q8o9XT6wRpk5m1yGAqe4G0zM2C+SR/IvoSV0qCH3/58Xs2BF
VVOfKszfM+jz4erbMuPF5OiYByTiJ5hK4IWRqo/k2P4ztFqOhWgOtcRoXMnIaLubfO5A7Ng3cXAG
OVvT856a+cIDuFxETGIR9a3/n4DcX6iVQ3vMxuqXgsfvl6H+FDRFf5/rpCZM3TBIAhk2QqZrIOlD
m9TEhqSCvZde2tls+G1jDIXD2AgdvpIrl+lr9OkienRfjQ/tjlBX4pJ1hrZR+XFapzCmbTmwXy5J
lxiPL6aQlGzdGUVlfzm6PU+7ApwrnS1d2Zh1OTzQsVLg5IKSFKWKGhoiNRIto7I5KzwfcvQzULLX
wgrEzc0wKtDtkJ+Vy4RJLjt9f6QXYIq99SutKkACvK4HZDUvu3DFT72xTcoWzqJCRqIcfxyhK8gT
veJJYc6NpPIufJzzFev8B+upu2PXcqRL6SW7++oTuYHYG0nxhgHpyIf2qy3fD3S18KkcyUFgeUpu
tssATRM9qJL90edRJRImCduGY5MQcYGMjc4SA6qvYfWl2xPdNCQ4P6bdHwMblrYdKzGDrO4dwvFY
5ka+++oGanr1fl/ZKKRkw1yJJA6yMa+v59HKPJ4b/L7WqyzJeJag4s33uVKl97NTzmPYF9Cd0nP8
Y9yb0zmaAPSfTmigQOX0rWdlH7MMBGV3lBkyWFvNCRfuoYYoAcQDzcxMLllYjw1przo8t2eAf594
uxpatHPJCU/mxEFR3BBGoXNdAL+7EO7aruQfBy5gLaTT7uDhMHk1In2ObZ4hFykp+gIdMSYZpDTV
exIqZvn1+SsiAbZmWNKEoOmmzITC6MlH3S3FU20mgTolPv4pALp/b5tmW2/zPGdE3zF5EamJdG+U
loR+afLjljdFIXep3D3cg323H//B8LjSzZekHZC8OVtoyBiNn/tWbZN5jdxdoIdSRxN/s2lFdXWE
2hT4ibAycPM4J8Dhr4Jrfzj2ITqQqHNABV/V9KCLT+JiH2RzAYxLmoB8N6bJNxkY4Q8jCqKO+tR/
hbFKGnYxr757ixYpPMPI/q/HRNIlQLX+z+jPY3muCIVyDLX6GKVfmwf07mm8jRe5mL6Ua4oubo1b
7Xj7II1HxGsJ7dhTgtJAivm2xyCpOKUrybIJYtFU7DyZdTGVMzwj0J0cPrquT4X1lFAxnLCADV2W
r5yc5uZxsBCQQVnP64PuKXVNSptQVRs9alybh6c53WPqCPeH4ioz87cMRBVQ9fVDmZyPAmNKLmiU
PnsWIBP2JN0xJ5ChzltG4qBDv+//s9l+U5CuiaLVbLeQNenuQrskLv/WceYMjqNtRb1Yls6Qc91e
3UzhzcsNiZUSITMW/N0FgTIhtxI/WUoffU0nKuIekR/lCMPJG2zzwvZn9AW/C1ZCLuYtBxxKqjLY
KE2c7bVzAqgSLfbiK25zwrPslO4avGCoYjbS9AO3YHxCZstVnAsFp9B5s3wSlrzD6I8mycE6Tf2H
EKJzPxxdlT+EVuzxQfEcJ7kpOycj8oDejtSU/UquEWnx/01cyVqewx/PPvL2jk+sthYG7+qjGobM
LYzcSOZ+5mOSv/rThkFP2W3Prj1dz4PlaMJVa6YHHDLrEJMYgr7iwnMb6f+50CGbuc4c6750z0Ka
baZW3vsWy5I0M14QDcYIIif1hLAcALwzZ0Fqt2ojF3WuHqhesuaPYlGJlu2Xu0u+pP3ITssIiOj4
iv1t4XufqKASS+6Zis299KzyOzw5DnzEXslpPivh1VKClO+D58jkUtEjpyM+hB1j30BfKM49R0i3
lh7IZ/6d5db6U55jD3cFW2AZGDUdCZ8OCtIIzpWGbbH2TdU2PpteBbooKPboJX5xNHo3wACTUi7q
fMCe+mlSFqma9J+/WnBO7GDUom1QL3ccpvHSCjlisa0ap3Z4yYjLOUOsb1nSsysomnqsL1RMiOxh
wt7h6V6doEX3D0MJdYLlo8tbNhV9UyiUjtEPq9p44dkf96i85djVBHyudza1iSk0iBwOgMNDdjAr
KoYzW1NqeFhV1kApv7YkgTWzPS8ZobLOygC61z2Fr9Ca+QLmMSx4duJJkqUARnLKMmRGa7ubd/aq
wSMGJZ/tmT9qejLkiWA2HvXZZSY5S4wc2p4kuwk9NLG73gtDkQq3JMN6WPaMHIFeWu2ehFkTLYeC
7HxaNmrSwQzTNwfu0VgC/BgtI3dvONcbZaurLu8zXJYfWrS3RH3F61jb1uEn4A1ca7rgNPbRWEYK
aldBG247PN6BYeHMZCzK/IuY7WNL1JYhAr1+UW4jH4hQFWFL1aFDKpqnVYwbtF3RnH4kbByTjGgP
+xaBeGrX3BMcZ2ZaOpwIiMOG6bjFjGZhS2TeJg/bidE6ifMOWEryfl450QgJOhQPypwJ//KM/bzR
TWOGczvt/eE+5Pf3cE5IQc91e7zGHAF7o3BgneH+DR1H1EE85uxcofyTxRnUNJf1SOkEffiNL1Eu
fzi/v7V4A+cxIVn2pi/l9rBUWsxQaGko/HSxRvMxaOXKCFnoLzCQc+i5MmP4bt835ad65szCiJwZ
lQJ20J2y5GjlvwR0TL8ADIZ6mLPk9uU2kY9Bigr/F9ruNXOgLa/tIO6yQeLgK5XLaPDK0+ZAM+bE
tCGN3YErLNHJqrPriYT7meeSyeq9GZ9MucgY8jAdDabv66BVjVG3OzxfrG2zPEIHto2w6WCT9RX0
JwCNftL7GKuh2nbqbaX/QYdIpXG7YNxdbWSv7/4h4ynpFPOou1YCQ+zkJkD5gXr9Jlz3nS7pwAnu
fzZ5oI/Ih7Pe92HIS6UDCwaPZC9wyrIG28KHI7Pi2Mzu5t0Qp+SH3TB/CjN2WAMxc2cWRqg1EnkC
HVsYpBsIUqz9U5kFMbKcV16zKWjVHn4myG9Dh2BnGBtwZixjLtFn9gMpdgn9K15jix9VEbSoS6gw
hAhRIQ8WVe1bszhC46eK4KfOv1oXrQkdXUytK3spyAOEdTpDNTdkMeEx8aXrLKQhDD6SqFD2/2zi
8EDU23bgpIOiYQBLGu4lFxryW43Jx+HQKCQ0vpJirbpJuMJP6e+B9rMcW+hIBqX4cKRIwcb+6BKc
GGxInQfzn67DnDxQtcD6/2Kg2lY6JHK0omcPmd0in6So20LZo3WV+0SneISbY2nEwAt/jtjYkZGn
+Z3FRLe1eQi9w8fpgv9Kk9LYeNHGOLP2qGN2ySmxAxZJsuvjad5itIS7CI6pMTcjhwepWUVrg5PN
kXT1YZxtFCcwTjHIXIotv8wUNtHmPqo4bKLjfeP6Miy3h+1UeuXgWv2xLGX0o5x6kuboo8VddZpG
7S3DO/F78FXu00NDK0/A+BWFkRIlGHtEzhCaix3LLwivSI2pzx8fa9VkUN0FyUOEen/CGFTSr0hF
fPOwObWj7ZsxdbRSTRPhNXmpl08qk/qBbngNdR960+AkrFcxWhaL7MZ8xVOO8NjQPYbBW69BkYhw
KRqYUWV1W+ieQ4e/CSQsqnjCwU7W+nR/21W9q5FQWP67OwHcd/+9Z7cjB5KpZIFwV9c2arWukN8E
HvZOdaILdI1e0qMGpceabZ5PuBufPSv1rt5bsxxsunZmhL5Al4DBWBG0Q5rbcaYmXPQPXnfkLt3d
8lgx1tmJ+cZmPsSAwjZFER/JFgTFXi/llI7/5uqqw6JBiGJVvNT86zAkkSEy9D9RnT/OgE91G7Ho
c36N9wrkOIe8CW+qEidue36CgLBffeZ010S1rsBKKW2FhMA/JNQdgcIK82QRx7HcwkZ635PxmR1r
3GBHCs+1uD6eSfCU9Jon2DVyg93wCvCTAEGtpK6Ry8xOqEGRXWY/y9qdjzxtud2P4n9BGaPe5N1a
kbIhYY/C7843UYt8wGeItNwx3tQqfXiVct/7yXpsO6Ec95IYi7KYROSv5ghWECGx6Kj7MFwYt3b1
cKqZXjzGfiSGbSJUY/yCX7LZkxaNMcFHQTtEdkakf4ESwGJ3Z7qy7v3nBgV2r9oUER49uti6uZyB
EgK4k/RNFaS8dg2fjnxB2/7soZ58+iChwp+wvmUqGUk0Olipoe6WXSYvOsqaSCXx5DrRjqWdqwu9
9KJf1Rqw5wBgajnFSgBnmj47ooQEzrmoK6q6elW0CfVPw2FwdItQ3QiIx3Lf/FKMY0Mk1sQhJc/N
GN1gsbU6yg8Kuskm1Jh5xsHb1za4jwzNvFK8rWbUqygmZHhdciHLmQRJA2IlLPeL6BzWGoAI+sWS
fxY7P+Jvgh5HF/gYvYiODb1/wqsx/hTDRu9TF8y/T2wmAWc5XaqXak18ZAsFpznAsAIOivLUfvQJ
BeyLnwR84HDKNNX88Fm6NhvwJ9RWPCy7NnVuuK+2bmNTYO/x2cLL0M8bZTXDRQcKTrBnR3HYSmnT
brAM7hv07Zl2Y/9MlFfaxVMnD2dOJlwuoMrSYQzL77cDCaTl5Av1fS8U8UtvjCDsGejRl8eaAw0a
VzOHGrVUfK7mt44isAyao9+SylUmSX3Oq+J++ybeDXN2NGHpbFMO56S8aB63eDC6JpsaV2IZp5KX
89oDEhDZP4XafevDqxFHqLv3iTtO+9gPRwq1AvG93Js1wDVZc7nUBK2ZmYbyomnWRW7xbYMiJww5
kjyqci8hzjR660w2VIlwp/cymgKx7TJTDWTKVZ+4YytkHZvzdtUSu2eCyxh2QLFLF45v7hXjBxpf
u1fgxmgu5YY+F/HAJVD2/PVZ/cghiRZ9SuKjGylh1hu5KKMzTFCwig58/VvMvz1IZUN7+Ra2NqO8
xKdKeWaTK/iAok/L2jtlldCpiih2oJXkBr+gHYdLJLJk1eEJXpGVwgI/gcPz12Y7Zl6PudPtyqTX
IldM/u/6uh0qXx91AltAUUnV/T1d1+k+TyP3QBqySQRdMtx5lM1VKVrGQKhF3nBEHoSXRNUI/LsA
t3Sv9R3YEQWIsN6jlFJAMzudXwMHsgIiYk/NkmXV7vY7oZCFlXSPCMETA31eJjkDN/hIHAIzjuPp
VGVMYbdNF4XAdcF/JKKUNstaf28QXWQOaahmOa+tcLTO+bWSMV6mmkhPq80sjl6Ziqfmx4RfD4FS
DehGTjQP/bkPY0c3xPfpD6OWMe/MoApAYj6AsLyQIldx/T7JQaB7nBUf4inHp2S/GV+tkHV4KLcl
tim1hLgSQzsCJslS4cML2ljAnWcygdHnY1mD0GOqO/8flLSvS2NGDhv2kse02wQKSI6dQuI37ZK5
2XI8Jh9hxx/PicP5PcmgaGq3VTo4FDb+3GCx4JYgFcU2UESF0h3DC8ZJpffyGfz6WnVIMx87eNAQ
8z+FEUh0FefmlYiHZ2sNOOoxdKpfGBxnVuFfkTpXVyevk8alC313j6rqDR4u8HW7OWRtRnK5Le1t
fOqeOOtmeVOdgJp/rCHid0MShDec7L3hq1En61vmuhVHJq32AtEkwbJnAprCHdIDFBGtKrV5P+2U
X29y8ENpkcn7csmqOByUhQcivIBJhtq0/G3ghrACndgJWdXUlE2bcwnwfj/iURU6JpeC9VKW7rVy
032/ihsKFAk0MYP8uU6AHzhKqKE0a/KEWk8FSl1M0EWWkAlOwWEsMf5K0JA7MHBJghgKRhojsUm4
CnEZJKWTF/iGOgznNT1VlK3lwXauxT60RKsqReE9JrYVAHHzBr2QCTYGkjqX1pmdimHZBytjKUd3
v0yJ68UL/m48SeglQ/UIFedBrpglAETvpmEBkgWWHXFvwzVGswFTNl+KFWwwNfVcVRK+dbvd7F2O
GSJ04dXiEoCRHawfl8PcRjuPf1SX6TsEYXDpFKVtjg0C6oAVyoAeP1tmqQdp5YJ28py4mfQ/ee1b
w4D1LthBeULl7K+z6DfG/iRqAwkE9uDrJ3LyfCXjqIRm40NtdF+gz1VP1ijmW3r5tNhqYHRHupeW
p9l/8QT3JfA/KYHFOG/fLGzbPpQeOySjRqloAR4fOgNosrRkoHykUz+h6hHVUczUAwh4u97+IgKq
zT8JeypfrVR3H7fOkxwEwG4MLoaJCaIJ+ZJ6xgdmp2H+XBoGKyeVtYLQfojJMo1FkO2fl5xs2Nci
t/W1W132d5aQ7Mom3ByOTmsRaDDzHukczLBWKnS8lXj5tiq2F0oPkZVJMrN6Sp2jLvKyFrMkj3iW
1C8OhYnXVaw9vmnogT0oRjtx5mS2Q9xeNRkjDNv5hQcVySiCbYnu0nb/edKvyo/5DudZ7L/Tdzcg
kAxWo3Rg74M+45nGazeFdi9g1kfOfZFCoXCePQy8S4cr/FS1OVwG/cCm7wmZ11k6UdmFjHdniow3
ibEmcLoC11tczeHnIZfXqGPSoPVC0But2MwoAzx0UQAX8ItzBkQkaBsStt04tDXs/qFkYG35ep0y
nvW2Xryx+il0YNOXTN8LhIW1twQ2oingVctjHXxcT96gRwiLAf7o2d05uV179RDVJRUp0Tt1LcRv
HGFA066slg3Ljwd7dPzGlFQEWzMnIOlGjGZUKGvx1Un1VEXr5iS2AGNhT/64BVwhD6aZy5JyKwXT
ps3HAHa5Q1E2NKl6fpEaWGGmvP/6Io9xjUqO463ZShPljzPDXN3CBtiJgLFY3tETnSWnbmtCfxkf
CpUEPEdrXUKDfV4L+FHIQBuCavzBvEYNLdL+KhgOzeYT5i+tF/vRyTn5+v9AtFVlDqdF1r2ccUkm
SIyRJwH2kRcDe9YNXf4gNcQ3qLg6d/Lc417tc3WaC7DbXngamu06FQh1JQ+sDMO6qrlHgrGzzyJX
VnwH/pXOuuiizAr6APt3cIozboXD8LEaoSt6qnKQIaauyMh7f/1AoXWDjt1trm7WWOgQ0SJYFZRO
ThfJjMKR6DfjsMG15hk0sVKcLpKkJtQMjtfVr2k5uhbAvXRMtJPbmof8VcH8pXB/ta+XSnjAQD1C
1y4CxxovOb7qTr2deXL/OToeAEK5PUOVRmGGQFFYtRbI1l3BnygpHur9FhwuJyT53HjAcbglDRZ1
GVLqvsw3nPmot8PuXD7C+rg+nOud5DUS+QeS/QT+gEYWzNn8Xv1noq36glycZclGVA02XK1VZwxf
a2wtUf7gUGMEV07+mBcvzRe2wxwcKiZfCzxwnSFviggwqo4hBkYEyV3+IlHuQpwke7a0+N2KzZ6y
EoTwC07l7o+gW8hY8Dl3dCyNnLm8uho6g3NwEvpvnJ/1rQLdHgNvliKlPZCNN2L6m6H2CohCEWEh
qLn61SMqlHdx2A4ViSIPUfUPUFyLB5UMaykY0OkF23D56JjeC+ZzNoYlptKY9RRxbGURqeElhhcI
wQaoVnmqVt5X85TMv7pJUDBTyNTy6Dq7c5jMplxyTCeruDtlNrxtmJOJ6/kcfIiCJ29mUhYT/yCj
iZkZhMXT04d/MaluorokgjbmVc/NXA6r7sqVRuuJ5NPOflmO1UsriGTmSjg8dY4Ki60Gigi5pn8V
z+lHZn0IHFOcOgqtYBu3oTamnqmqXgLIu0hLkH5CErpZsZuCcFbGsRQWznmL95wv3bHmeeptte7v
o+CPOoDrnP+5XcmM49gwxOv3KF0elkUWCvyJANcaIKWAkFBwNOZgETDNkgus55HEjVlM2C0OwddC
WI5DNuOWoDgM/+UXio4Qtqo3AeURIQqxB0xiHF6ICPYjD+mROZfADAuJW2MQACjuSzWuHj1Oe6I3
LzqkrLslWCVMw3FwYZKD5fDJO2eL1IkDfa+P6MbCOvSz9L4Ct1rjsYjeYbQ8dlzfqqXqO9Xe3dA+
mzsxcNBREzR6jLLyoDw6RszZ6MC6NjJs3YbrqbwyvGmlXVwqA7TNvcKCCs6y3ks0/s7CLZnhtF0Y
aJ3ldlkmPynmz5Vs4X5J3izjpcvwAHCQxIGyrTd0ZypE6PGtamkEFvZBvmv8KWmb0/QxILrMolM3
xmOLzfVgKRNWWLqDg72oBWK43qaVTiqoNDrLCF7PVU5Ct9DUVzCtsWHpmQnPes5aXUTyjvAqzJ0t
bAY+zzJ0v6kY77qhODRp2MbMn9X5okC4k8dbxbkQdeJQGQ4Nk9tPRQVZUCQKK0KM08SRyObS+Ftz
litvig47f0FqCkx5Osh3vnPNRB/pj/1ODYHkz8mtOMxxJ07QIPzZaVJlVuECXBrxLn2IVPdJl/vm
PRji3h+5/3nvUJcERCYZbwwN7rQLGslomtU/5GI2Ep6TUeCwDKC9BhsINxprpop4dOg8ILVN+kQV
T+oT4OI5e3rObpOQ3sOH1xuM4n9vTwd3iDY2erO7D3njVPJQs8E7KTtQunwWDsqB5VEADkNNFjGc
WZ9bG4HaiqHQUCLsfTl8NTo8qLtXwMsgi37xehy01gruflyP9qMknrIBiHEGRjNg+xO57f3mFuDN
jtNmyj2Xhiy5GzxIACJn2oMcqEw94ppNygHiYxLjktcBcTLhtWta9ZgLE2ScXTPdP9+iH2azYLyD
tTYGilxhbj04X5xG+nTPYo67dVwS3p6oB0VFfbSoxoM122KDjX26k3CFRgm91MjsuUWKdRYkLEPg
PXajzO+d80AK4B4tDKN02BwyI9p9gVStDt5206WDs9wsWTOCfO60C2D/Tmz9VgkjXHlWjIihLukX
vgQHv/QQhvGr63d0AB9YMnwN+vQfgpN8h4WXDEWlMdpqqH6i2d8TZVeRkj91+MLnMV45Q9DljuVq
UkyLxbCBfQYYnRYhEWWWcFJKKpv6NfnFY2+Vj93O6zD5MbdSDQet8ytvxD0kt5IMbBHmsDAflv+q
XGM+kw6tden3H7NEW0kqTAG15HcQnEpIh0zX9V176roTYNgZ98schlTxsPZZceQPhxOrtu8wnXuF
WkYPxlMLVUfDl8cO1ndguEkna9karWyoMrCtpATMnFEkrbY0VWHPgOLhuVE6iB3UzHxDVPuRnOJb
qPiK3Jc0Cc8mzZq63TUFIOWfQdaDg35SvklqtCeHdm+ChnQ2JosaJgPxFPN2GTT+ZjeJKNMJEdlm
iGsrC3Wr7TSPIRZmNSVps8VcZgW/RzU4RKdFifQFX1D3isesebEifKivqh0ZGygji/iSczifnmXn
aukVYCMJOhEYUQFv2o/kjVe8aWIqcKdcmA9CCXFjYrhHUAgwMVBwAL6d6GtztqjHOVjQSfL13Jv2
W1UIK1ZOluiRA9bxoq7MqmaxXED1iiQx++1m8LmygkfiZZHddmw5xnNiIzrsjTYjxGr1rJmeFd+2
mxbukc3vBjzbcgFnBaW4jZbEryRHjsczLXWct2MiMySFmA6y6ycpPUxU9ywk+kha0ezNCWlKjrxk
eUFS5bel1sWGCviSIn9paMopzUWMK0VqptfMFmsWXxzpgi9jK8uMsXNUiSNVxuRyHlGNc2jEPc/s
PrMaCqTSEYtJQZ3pYLXnMRW09G2G6AtnJGuxa32UeHvWfX9OvLh2wIMZx738IojTqIYKpCBNZ5J0
IQ2sPUtK7ur61cu7w5mnKvbrt6vm+UhKjkDpW9Ki7oCj5XpS9CKZo0E3P0Tu2Kh07Q9pq8EuIsMz
8/fS0yfuiqgxS0GWYfAHfYM6Z5e/vRePY8Ldy7oC2lxm6+3kuRzJdxMEyV1wv9q8B+76VbI9t8bc
ejzTnoP6JnPxInkXWXtlcVwLXbg7WKYP1fIXviW2v000eRQZHEi7zmfvVuaRzicJWq+bN0ZKdMds
l7exQ6wzxDaYtne5TPJjt/F2PhW69AEtwZUHJWs0odvYXgev0978aGcq/YV+DUfbVshp+73k7sUZ
D/86GZ2R44fe4A5F5Wp9lIA/Uh8l7yj6ijjq0nZapr+oXUMUCzPquqnolWfuL3b5JwV1q+0/YYb1
paiNay5yCunxJ1ujVJ5/vPRFOLptNPfFOEAOLjnBUDeYYY5fif7feSeWx1uUc8uvOKDAV7Fd7AkD
frd09/6D19S5bmROM/OlYLLergUhp+oCv/aC9CEAKUbwPwt1tpj8l045c7RpzeVEITmqvQ1Zptmz
3HPiyWJFXlLZpJ6rF5htz5bQaSWKnJMCRtkNOLNFBFh24GY4tIpI9KD40A/mCyu8sZHg8w8QGl0u
/OcNBwIA6pgoXek7D5Xp22u1lKQQdk3S24N45forPDca1dKPpSS7hyAkud4+ZkZJRHGhglJuQiV+
upRxmB4UoPrvE1GRgN46srZ6VEt1/Uu1ri16Kk1/qZrmDO7jdJspi72ADKEHYEkWWJGnxgBRnWvS
qty2s3CEpCzYZ399iY0vU/zxcSAVJbDRU9cH50FJ8D0D0g2uWqJK3jaCu8SrXBa1oaUnLeqXRxbj
6g9A/LuzXxCIG+4ySyyEK/BK6OO0vtYkBYmriX3SdU9vY2kMxvOIzA/hCdC4NKPxFiRmI6dTh7+P
JQI09MqPYHc/E6TU7rdMSn/aQIfr4wQizLYQ2fLlPFNPdfgVbietXuYxIPEG5Wn8ie28t3wOsFnl
KE8/1bRDFQVB0qaWtFsTfwPurtS6uoCRF37xRVkGjdc/7Kc012eo5W6VX0tlXiLwOGjJ99oH1bNr
7FOi0bOHCatBKrPvDczQWYFOzekNJIwnyHToJ2i+N7YQRn4AAF89a0aunK2JvgNsIQOICrdwyVoP
ZbTtvzWzOKbwa3gvMjCU58v8MmivqFomtFlDOsHHj+V2WK9B4Ei/6gXzuSHlN9uAErBgBlsWaE0R
tFuC5YJrNGMyoiZreeLuT2xelCcIGjMbkgIe0ggCJ9vucC1V1YJiwdKc3xR20KH6PJQx3poFv+gS
xt2FxQ8KMX+aD5w3QtOHGtY9WJin/JmklAjiUyVU5ssP80R0uPGqFvH01l4shYUp2oiBceefN7gu
4a4rR/6LlOQ5J9Nrsxk4/iuleeoTVBJcJQb/AF7R0U3e4t9d+MD1CPVr7WAZnhnX+a53ntQOI686
MLyQBoAqB1VdcwukAivwinOJtyOIwh9NgVtztt07/myWawA1cgdBNZOS2+0PILGCmfPezr6UuYwA
Ijp/JQU1/tsQZJxhJyDbWeteqdixT/TMHQqBMCTUi3sP+G0Wg8j9HKlX1fE4CUZZvkNcB47QpI1/
bdX9aWBGKOjZ7btcAwp++2/t6r/vkmHxzbGC2u0LUb99gA8WUvmPcQmqOUQ1bXpz0VdAZpY69hce
WrpTXW3v8Ri55TNjgRdIxlc8NsS0oqRcLTLq+pfCaaRNPJMGPItWHUn5zZdZbHmILkAiH3WwTFBE
fiwqhHxSlX1LsNS5xy3kMBEIIXH6SMZ17VI6jRhSb8GJXyfTovU8hUXBn6+affhF/Nd8dqE9rUmD
cvZ4paPhR8e0x/+MHtLN//wRzhn41dN/78ly9xENIi2iLNtefhTOKz2uowUBrgybZ5ltJY2yY6Ex
E+d8qa16KUc7CMFD1SX4bFJ2bG32+P75vBHzS9p+wcnD4zocY4lCFREdkTqFBztVLVkK8SCiAE7h
hQ6Bc39BVKARGP1ge2CAsUiyuCrg7OGbqbHfa7RDMhm6b2yZjntoY1AWLFIfzUqo19Ir1vzkYV9D
4or+lT9msL2ymgvAB6VOWJ0ODlrjouA+qA5UX7Gk76jRA/J9aqpmUNY6y9JhMiNMd0S1jIxjYvLI
IcQ7EGv0QQDsYn56YSSL/FHIxhwLkaJWIvymfFbyZoLvSewtDrRd45QKar8og/zqo7fbpWeE9AHH
wnq1idErT6Dh2uhyc0Syvy+Vsw+dXeHhmVfG7wjFveorteH46KntHofwyjHvVlxWiypAU1K5lshp
HwLkcALL5/blbj0ZwZw22n5b/HYihJueZJlVO+Ax1sqVy88K/+taUFqQSVcz1ImPNL+SDJIaxLfJ
jZwFUpnK6LFgilr3Lu2W11WjQCmmAtI+W5So2s4wR1MSHwL7yoysrSl9z7Q7w1JIu9m5oqlxj2nO
TmD+bfjtDXLbAijwVXeIEBFo51kR2H+b1KKaS9MNk4/DVbp9XCIPYCIjgO0F2LJWIBCTamtybdHX
ZCMPxDZaOAcLRKfwl9/+hMFeJJf4z2SZ77eCHvX2ZhCxP2JwsmfPtO07U39QKrcB/kCAL2SD5bFZ
JkdaW6tp6DTDD618AZzkyjw5WXHSa6GRLdlQYYhsiAHQRk2iq7rKGWeiYuwKiiUfiIernbxSKymt
vgoloViArhzU5LtQmzh7Q2YEgVixE42BeHEmVhu+FqC/mmg7qzkBa5ULNBMD5wrdS8hAraduW3MA
rOg3pel5goAv0/iq1zA6sG9C88JQ6zev2yYG/Mudg38IgyzrsbuuYoiwC5rYSEUa6XA2jTKE9lAD
K9FbbvXfwqEmyX0QqOPpWXq+hRdVHUwdRgGvDlR6p6Pxvs/lZHEaRxKcWN+4n0KcoWfSMGP9h8Fd
jGzaETEVUurb0c6++ftNRaPCffT/GPLFHQYshDqtH7A8nNiYKIBbvfB5QKyxxRzTioD6i6ehV+E2
G+TrI7EmnKRUB6XA5fe/NxWBkoA0R8eEghcw6qVZev1DRrr9WFca8NvMngdpsVdbYIK5Qn92K4iO
OtLCl/+4LMHWfZCD+zIfBr0FAxMAuhjCdgzi6IfJlfQy5NKm9rfYHFC5CQ2h8PpNZBDHNAaVUf2k
YDvKRJoGKeIRzBH1g5xhjdFbbrjAKt9Nb1hOCq/mozx5DWnBhV+foLMiGIK3hCKuNWDuqbGDP2pu
rqgZdoDHIFnmBZnwEo/Gu0RQLVjhHJWSB4hqp7+H//tGQUDyDPZtK3d54I24dwkgTQcvN6MT84Mr
OGPXxP5rSvify1TvF0IFvzdlCUcuRKq1ms/bPMGfCzyjaIspGkr1cJglfJepX9DzNYTU6QTNQjts
ERaARnwolB6HOQ/BlPXkbjfiRv7go/1kMfq/bGnnN+UhgdPmScJ92B6mbYKUR0//FKo7tAqIXxNS
ly9iUjQYwNS4UdGmTv122NaLWx+WadDz7RJ5g4r7kzPZLQDI98GP2iNe3/FtpQIYed9sgYfrc9wu
Aamknav6+ZaJlxkwV/hbUKVnuZLgTteOi59ClcQOie8pJHj+4HLIJh8l4dhm9jIPSaLSNIs3Nx7m
JoeqMHrZa8Edu+ROpqpNpumum6VP2cCYuCju1Zer94V6GAwbv4HLuC65hV554q2UR+/5h0OkO3Xd
XI+1Tv0idUtKkUjbWrlzByzF2qlZ8syu7Ncu30i4znyeQKAa4lGWsVIrhR3XoHFPIjybj9fajfDN
/BaM3d8sMYk93pxiPXzvU+wo3c8/eObAoZSei3OhQItUHS/YXMhXUzoOja07fGUkzw20x80kQtxv
KRuTCzpEVIdpXHBQwohZllIEgFfUmw/GSmJ0PdvkY1bvbdTFPjg1JCvdL4igLnpi7Ep/qdzo7QrJ
Ifd5eMu5oh1y4jgjE3M8ohLatgKxuKmZ7YpRM7kZcU1m482xt86WbPrHZXbCex2hvWAFF1RiO63V
a+z9TmvqN5X9byHy72tsDYzrfANi6F/BqhOTuSVwiQ5bCndT5mccZsQfC3ULsFzHZQM5/sXE8g75
naqQL2qHu3ov7ZWNIeeqVIo62nCeypCB/NWiyi20XWiSizzwOvh01UTj5GMafyr3pWrcJSpFoyyp
gWCKyNmULGiTpGsjzlC0f5uIDa6Gyxwn/+zGJ8g9JNiuRHw6ndjnRYcCzIqvR2BI3UcOg501hjsa
pnOXpIs/JfvVw8Bnx0C4nFUV2/ELU7fMMXhmgW5voVS4rkvuMkXVu3NV0lSsIswPac0l8r3/X7Mo
AIQqmDJ8Rll2Gb6DtFNrhIc9OlxOlbWmoYeoIcALHk7WHbCGfl8Hx3UcMxIesvJgSDmR8HBYdijk
BT3FkEtfAaat3X6hfdNJsWY9FTKWbzCTJpFLA95sy7Y5USN98kLwuY+Z572xh8GUuxx3Y71hjeTK
B8teUWELtasy32IsD1/vyS74MRduSjrtteYMvtc6qb8EYUiiPTqSfK7OKktcuUJh8Zx8ExByB0L0
q27WpjwGIp23l6qnVrJ1nR9oEfd7MtAGw59IdxZLhRqXiRED7I9Lq7B5BmBVZARysUdNDVNjywvA
LODBTAl/6nEcZ4tAiel9IeXBnfTpuCIIrMtmXINO6cttvKY0Vy0TgA0OTw81E2lmdSW/ZKNu4yPQ
gWRvh6itCdXJTZNFKbLhjPgV3jFGiqqXDPCO6znaY2L58OqlGFLiHOas7xsQYiIsX37BKoxhoovd
fcaxmd7ekIOhiyPl9fygwi15gzKNjEC3rPrLNXPPaD+Vy85zgeGrF2eA4zbcY34U4BJo8hNiFP7R
3UXr3XfuxdHFE6QgaOaqszSm4nbphIKXCtGctpBgTfzIXYkfLgCdBXUpKYjbJX/8u/a3ob+IHj+C
q8LdNsJdzu26N0k/3BmSHhe197rt7F89InUidPN3Yvag9YLX6g/DOmYCE6LzcWIyZI6bgGUB/HEY
zvd09BXVRbgTdY97ZKj4Ycu9F4ZX6nsesefwuDPPbD1N1NYGz0yFkdbSzCc2f+pKEJWCHofB8yTn
H2DCxz1/80J1SG2+rugG2JetdprzNDudMLnj+hA6LFDuL3PIZ7Cf9NKFA8nxWBUwD498UbwWp59k
Rxe8H6JMyWjwxREPguUmfgDcG88j80god5Hs8G5r7FIV2HTQQD+Q79ExvbW6veXHA7u3kXzpJBWY
mJftX0m9J9tbKvv6dnLzBNtKiQTm7vJQs7yWWjdtczAxXYFvWy9CYu3d5NBB/awe5ZF1SDUp0erX
S1XZOOCnaC2qkqItAD9Do2btAAZ7c2m15fvuLivUOzF2a4sGBU6CXGaEJ7qhiCoeLVIk+T1xpoM6
SVb3KLnMHGRke/ykFI4XM77NCoNYlreXNW1FUPMLj0EEbZU+5KvqrypW7gLrwi/ZYuBgdXey1mMz
92mhwGTqyYamW8Vp0m7lwRc7QtKhusWwipgv80gwRwiMzj3210Kz4lmBFGxQ5kSG2+ms0bObXe8g
o5kb7UhWigAb1HFl5w0kciwvG0hhMWwryxRw4mDZggty3EJbD82aC4C5bEus1+MA1QufYFtB5nkw
7KVkj3bfMFcUR+hwVl9YTfEDVv76R2Yg06CbmZWxKYfzeMpx0hP5N+RYgf2ycVHyteAWICIdLGmB
QJtNudDYmmHFNTw7stpabK6u2E7kf27v38XWrmMBLZ4hg0PMxWUozufc6rnu+7EVxR8xa9L4fV9P
GbrVXdP+5mW2XOeN+EgjWZ7S5UKchnzm2hUHyl23KY5SeMho277OVTz/051xeMVEboR+4X4LQXvV
xczYKYIjkCLZQMmIIsmeXpb9t/hjBFwSwPG06/2rzd0jfUnZDgRJJPkENXAQ8RzYoWxf4rFA+nEO
/i+ihsUMPd/M26WKiC38Hj76NQXPP5YZMnzuMpoMnjG9ic8Z9G41eOUbHBJglaPgpBlyU89Kh4uv
LL/VzquGI5SlBNTKFx5qbXqDxxiftu2gVwPEGsq7mQ00iorApOMuoKVrb3jl1BGN8hVkzlS+rASA
RuRWn2l7aAQcpBZOHfCkopvN+6rdhMSp4yA8pIoxH53XPpP8yS0hhLa/DAzsRq2PMRkZPq/PqYNE
cWZwrR8eX6JwdE4Cw/0YF+SQhexUjU2Us8p+RWXNBygPMX23PAdBUPMueoqJ8tLnrRJIQ6Ynbz28
mq0iiBsyo2SCqrFGdJvR+AQ6cr96/R0fIyyYm2pOuvBSETEaUPyMwNAq65RuH8zQ9MxDYAbKs5WI
xYNA8jr3cB7ZW/cCV2Q6LnFXdMaVEg9381R6oep06uBztpFL3aQ93T3ceJWxgiracFaWgkkfHoio
2I5cpI4Jg0VtwcKRu3CVuVNpBuhEBnQtmEnCAwCpo/hMIuhEQL4gfMtpJwIWjz1JmbTOEQrmWnkB
JVWd9392wPQoJWao8JnUy9Yk9CrGwVsZvQcz8oqC7aVOduUKD1ILugGF4y/HR6Qfm2Jua1scHwjr
8h2BaaqSOhoU7ESzlYsKNrPEagCbyiU5Ci84mTK4kJl+umZhToA5TuQv0nK/jXMuGfycg1FPWpyN
s+UvFA2sbSzFgGvACtVt/dJHivVM+7D0ouPrQx/wbF4ShXhbw0yl45T5Q37JI9l3gHNQyM/+06rI
Gf/TNezlDFnHK9Oweg+h1c4P4e7ZY+GjdXjS6jJCwXk4nGHQvv8CarEe7L6tXLgaHBYq876gMWtX
dJIkh+2+DGgVYI0Rxq3msqGCzXUdARXWHypI3ZADe0yQyJSvv5aDGUwnW7c8m02sJGl9Dfk93wUk
buJNzSWcu2Blbxygbp0aqGJ/1RrWF2VTIQAA2bcrz2Gk2p3gviTWR2QN46BUTWgLh2gqj6RqXRnh
jqfkmCAAb6RF9K6fD8IKLws5Fisee1M8htj/5A482JUFqIu2+ErBXOhTcC56RcQtJV9iS1KE1WLb
D3Tf3vcRu00Q8TdcXDBl76BIQVh1LyZgCHv7VUteD2V67+Ty4m8g/2MvbWAnJNONOK5T3ASk4lch
/dSnpZFGSe1qUGmB9LugyXEREAumFG0RHwE/stziJKmelaJfzBI9KfqtG5c4I1e5FYhh3gZ7p82P
5+m3gQRhGeWIGPy663s4Ze6MlquMX6k8miRxqnrrMwGJnvlL0mvtkqjryHIolyH6qn+EOSulzDvO
eFMQ+/vZy75Xr3o+JZBdVbjP7zwrqjDZJY+tKpOxBuPvLAg/+q7dW7RfqnSzG4IAvnxRbUwsVkkX
KZF4crRejw5zQCtrIq5No0sNoj3xa1x1JixhlpNRdh80RRSk3BV81CWKX1FkBsqTbpazas2yKdTq
0PprsJUUhFA1qDmxrwrJFHzEaELsbsSgLkEJVI4EZnkM+sHuBG+/PpNv2mV6qu/ekUlQzDV9Bgpw
FGlRaF+HBYdXKkp83SUJCuxRl/S4Z97qb5VUJ+qP3k/Aj7SokIwdCyPEjO+Pu60GC9Db1ZbgwODZ
9aHKKJW4BaCWne0SjM/JuOr+KK1QnSA5xZ00top3nSzmOLW4E1Gh8aOeB+X1yP5RpgmykENM0qQr
rp0/kpgsWq5wlh/QUTWxgKP+TxXAhb7jyqqaNuo7uxOVlxEciCDS9pqCWhEfJMRHylglDaFvYcKU
U6AW3C5m56XV2snIRw1oSKAlHRFWOgfw0m/r2djPkYJ8XTjYR1rmGXPzS/lKwTB/Rt3cRNNUR1ni
uBV486f6VsPrmi5TYGhzTfmh7QJk6i33SHWfzHdM/JKrnK+7VQ16xk06mFQ7355zVmFFOdWdHfE9
+pA+WMV738asZgk51BTdZpCBwIHw5/oky2nhzagmCKNHSoMGmUql0f9zgLi12onIF2X4RZQRhcDW
H8LhB5budJlUoGR7axDZgHzUQcWMqw444kpMsGe0Qb5V+yidD+o56g3Y/yp/b62h8GTyvPXKaB2G
75VINE2f6YEsYbx2k5mf1J6dLMhNYHEV3WJhQzeMTKPDiM90c3LJxgxUjCY05RpEa2va5jNYay7t
mzIEMkP8SJzT364lurZeEc5X5pzuettym5K36DG9Ascst+9uhNHx7Awwb7d1dQZwsKp9qxpInrtZ
xRbPsmIJN6nMPLZ/XZBDpbADp2ocTyaDN3I9UmF0Rafo1ZXjZotlhUbMw5lP0WQTRsFfCwTbZ35m
DWjI7BSCsqmW9INvKhP3TexxdReHZ7YeJeG4EarhaAmuavFnClxQSX9jDxPjtVxjRvSHqX+D1A/m
cy7ZT6dI/Hg9rS06EWlNCm9h5bCXTdUeS8YePjVPdve3J9WgLoNY9WhOlf3BpHUJu84lbYPx/klO
QxLi1rsm2DuX0J67X46P9KgFiUjOmt4wSgFVv8TBM6tGw2APofs+Jwct1bgfKAaOR4pGp1e7+e6F
qpqUtQmuBNVffoOA2/tj8XjpmEYYnwSOXP1zIBm9/1CF/l6vY8+lGvy2qBhGPtomJO0i+oCEL1u/
obAgjZMBYmrhcBafJ200/AiE33a0DJNPlRpyBKxxUDLknNdiT/gHpIeg14nuDxmgzRtPMjGsgSsh
IQ2NLn1u2y+i6fjXJwUDpAWtKHBd+2JsVU9ZuU9ULOiKwy/7P7gLe1XCQmwKQRXeMFyDF4YYhvUw
WAcw8gFS7/Zr2xHMk/ZupbXwFNA9lQJpowz7bOYhO2pz+350586ZP8ku+J+zqbe3/I03qJy57Wy+
aBJ0hkownFbu9Bkw/3w4SqY7JHsKrcFXiJavN0j6ekTQL4J8OpTrqnM/c/Gx6DXLkt/4vHaCCzf7
LfjdA42QmLyI1VB1/Fy6q8AXKszuHtxZ0jH7N+VLH5waktIjJUuePxGZ2KlVT5Nte7mi5EVuvNXn
b+QgPDnPNe42FDDjFuGLgeuaUYTjV4XsZpfxq1viWwsburwMBXvysI1C8h1kWWHfV9sbhVonnthv
Y9aTv8/hXkcthksa50k1B7y9fOt9hYN9BO3IZ56Y8+jBZtlQkPp7F/Bqx0Fhcrna0ZGyP6pZexiy
BwN+UtGjdXPRVmTB+9tpgwovDQnAROHtgu76twohYKYWl4tUUvz7oQplufo9nKETGRYHAo2k+vRM
3YJidO5a2WMDXpy6a7Nu+e3nX24eOdv33ZUGJNHbZzdvG7VTf1REOrnWGZR03qNDFI50Sz13w8KB
sD/DSObBOwnr+waVRtjVw3laAuKRyRaojVW4jLCEHKFqkFK4xxMW9n0Irh2cyulSb5H1XvuvAjLc
CnIe6kyeECoCO9m4ZYZUNGgBuJ0S8hXlx/me93lgNaMUAbeFnCjWP/GNCzQJ3nNheLsoDvI/MLHb
BxaoGbjenjjI4o91N7mPYGOjnMRWlS3adO4gvbfiw8NuAxwMC4RbHp6v/DDoXzxdKLfFacqwkae8
p6WQLocjml1pAi17x0IXtEs9BUh9ln/Tjk4vgnpC/OprBFzzR8BKDb0qbDVbLJOrNKc1+FgozYuu
ktpN7gvc2YQwoqzZ0t8XwF/Sq2wiU0IHu95Yfq/4wtr16aV14lxYuuUQIscRmICY1nsSKqTokJR2
rkkJ7XaH3QdqSkuPJkKK6nc9vFdUtgVXL6SX8C8Zfn+S9cA41A5v28qZXehyd5MJyodKjYCViToa
jw9Kuq0CW8xpeiTwA2lPziSzsjAlBV0fI/osxE2/bRJDUzJQ68pWk+60XkhK8K5GJj1qWjcWReiX
va19kp3MxxvhPeTmkN6R9rXY+supFXWhsU54fDAQx2ZnM+aadWa3q7PlVRe6Oat47b8KQ4ia1BNE
Q+4eiUYCsRoh2sluiAONGsYy8VD1TRGJzt7PNUe9f8g2CSVTD/CjL5dDzCuopYOZZpgiDI3ueHAE
wL7FNuWID21MFGMRMUUb+iA7J7qgfl2/NVjJ4p5tJMW5uV2brD8Z50x4XXtXRxfFJlCAfYgFF9n8
vFDjRMWaO+/9ipl4slHxHTmvjOv1osgGhkyuUS3W65qnBg3y/8NcYBaiA0SXrqB+1lziHy8k9U0U
7VuNVXRFvMRS70Y8vjRk4p5oUHIvgZ9pflffCCeCj47X3LnApi9EJSWTAoTntyPZqU48ZDrppQv6
IpdYvt4BcTTsYwLxYf3yDsJEYqABWqHiIQa6eoEF/YUX9pjxZlMVfvH52sZ4mHGVZVboswv+gCw+
r21BOfXIQA2rrYjNSWFaeSrQob744EVBCsEZc1H6q5/oI5xarF1+P9/Mtftxm6KSqH1gAYSy1iy6
b4SeCMJY+LI4NxkA9pNOBH741ngsQwEeQjXK4o/WM8GD/SFxV93R0BrpKE/QSB7EWFiZEpR67eIE
qN+5gkc0WcnFWta4kt4XPrfrahZO0UF6VmfgPpF0PZ7APh9NpfgUiy6Rq6YKsZO6uIjNSCaWRbAR
zgKEC51VqGqHC2sMpE5ZACPxBvVhVvo0+EX0+OnO6ZZOnKQJG1KnEsXuaj/ssJrpwHAGaB4DnVEq
i2BmxdRxIJPERY/mocrVFXhHrVZjghTMHUsug1OiWIDTDzL5G5bqMN3yCL4ML1xr7pksPpPB0VS8
26ZBTDWjxBV1lfdaGUYKa/UQd+Ye5WG3JDpq+0qmFiPde5TlJzIFCnQIQ+5lPA7q2PXyJ6T0P8k+
xGw7X8J8iJqi1rWpNaiBq213VEIrNKwOORO8UYaI/vjFXzsrrJPp4yUCDwUu9cb5Chu9+O3lKyP5
DZFZRSM+80MTFrxQCNFGwkvUgo5JEv8EisDPaDFGm+f6WtL6srB/p3m5MA40F0Ci4fOmlHMy56sL
tij3pmW6K4jKkie91ctzyV0YVbEywdbKd+YtEW+LgtLZcOa2Krsw1VFKSj4voqEmIxyS+ug9EdAD
n46nm7dKzp53aKfgTEAb/+lkvP4rPDn8hpWYdfpQASX23+m6/WMrLwiIX5IkwWeXsPAoBmRiL6YA
PBl+z6LcDxiEksLNab3VuGyn93kbE3aYAfZ9H8391fJhnW7qIS5cD9lKtqxw4fg7Ygc0oG4dr0ef
D9AuKa+O0M8xmoHEPTuCtBo5e/G3Wq9L4FLWL/8uMGRLIr+8OxPVOneh311PnEVmA/9PmJMNk3MS
PNYpglDxkLZA+vxL7+ZePG2fDpntGjMAWtYW8nzMWAIH63gRRL2m6k5x3ySq//YpoB1ANVq6if85
gMT/pRFzVY9dXYqprtJUQkcad2ggB16m/tqYQH8GnDDjnvRbXyq9+M3SBOyDLpE8eg2fdv8sZ+tm
aSCD/AgbKVQ6QZEqJtGW48DZWzUZdixpVU1WJvMaiMvphww6fktIVOoc4lSSW3JKtrP/mRgK54Kh
oQt11BKajAp9zGI2Mb1kwCuMMFRRrnFJtjl3J+8cbavQQtt4+kWaGbnqjVVMhu+p2VX1Na7c6gKS
i1PjzOqLkXp+Gpcg2CbBar5DnCPZYA1hPEGXl6lgQ4GfJVl9lax5abt6WZtOA/NUgmtTthlRPMy2
yHaaRXUGPOmSmqsYlexODYMkPM626YthV+N0PCQqFB/sg1z6oa6noyE2CjDpYWq1UUYcKtkfxMxX
eA48UxmohMGhEki9YNM9wD9UeOMH5tqpC59M+FKSDgEedbbu80jj541Cg//0wQJHbMtDyw9yA/Fb
ttZNn9FMgimn4nytLIlmxR6FoiH1QfZVS3iZIOGCN603kdkIdXOBW1kW5D3qlYJlr5GoeeDHtDMr
SOmmXOBgF3yrKk++CYis8A88dlMRUhMuKtxD/R3VhcroUyafjGy4pV1DXfYw8+5FeR/V3JUxchqO
NQqBODdPCFzpVNhNaytaFB0KzrythLk4pjm53XGceWzkvCdM0WjWtj9ucSBa6vVeYWw3BvM5PpqL
fxEqZwEHTH0TsXZJZkwsLgvP6r42Uqez9ZNK2OpgqVPTrzuWz2zuS313MNc4mfgekfNUxKdhvTFB
OFDqk/VsuUlxddTKcztBdi1oUcLthhT8ZiVIlcKsuYymfv9QD23azz++MD9fAaLZwF3EbznkDwOo
qZ9lK37aIGHPnta3hKSNxr+DfrtjbwEAvAHWKAIlgJWwr8U3c6yylMW01DsIgppHkiyKcUKVH1vL
nRfuasHEQKoKgjBnpiJvafXCs5do8NepHzgLZ5JZWJbd+8B7ioAFodJcR9hrm9NcdJYZG7oY5tX8
b+4lrtHS7/Cq13ZtaoNyZy/2BzZKwke1cTs5uMu6z1GsfqXOojktOAFndAg/8+kQ5zrprY+BNwKc
pVIRTaT9bjUfEGAi/+1+VUnthE4sIwIR0KME8NOaGYS+2gSqerESM5uxLqaGPyAwisujZE/8dTBx
sJ5Kdm3BWZsHR3lnERUXcSxg+YxtE1SbtTE4ZFtOUKzg+yrrRDTOTeORPpK3wXpRAlHjDgBGzVoP
mxmQFBpOU5r65hsmEgsLKJ6Y/Fj0mwAg8iDTl7jjjbB5wF2vFUtRXLFwvyMSmwfnFGERQtvGar2d
30Y14YJzM1o9r1nF62ZziWpy8s+qJ0Av4VCxZXFwiTTfIe3T5nsM5j+nUju/qggrsinzLPRAw8GP
ABcIdqSyhpNlnZ/RqB8u9YVMQ+rUBbsmXR3FmrBn6xfUUrdMPpCoT2uPqS9ifUSNUo8GM3QeXLM9
SyQb1fPrHgxFjyHFM0wJAA7lSAwyj9pI/KdIrB8jTPfSithKincUT33LyJBojr0JfkO0ZjjApe/z
2O/Ul8piwXyM+oCss2HBF+H9en7cPsOsKjpLF0iDblZj6avr9kBnk09abun8pjN0b+K73u/+5A31
BMIDXhy7HL9pZuG9UgE6qoDNjUKwFSs0+uIu4hKd0tNuXwK+E6Uo3YD30jCF6cJ3zksEkJ2y7JUf
ebkhMf0M5yVBGLb6TCNi5WMh2Tgr4PB4LLc8D89I110Q0BTkGghO8AmydCRHFtbtNx3snvef/hCb
N+I1F3zRvyI8J8EDr/RhVikk3KxlduzTQETsC33UEeubUuG99PoH/K4ClzDVdMih3lop8jUBEGbg
RQWt0kT4SY0T7SAh5RjacM585yxer4qgjVOIf/sEiZKPCkTXUKWhg9bLQJtpOHii3/BRoZxrWizf
RLR0sngBjUylwmlePkhUHxh6jyycYIPjsHSuQm4An753IKsXEPFnWgR5/9Ja23I3NmddpgE8zKRD
e72t+G0TOG9bFGi1uEhvtBLFgprRM5xRDDHPiGVS5lORi7QP/E4osnC0zmzRDKmgujWpUSsbcuoq
4gUjRmxWw4/hrjdh3JLOOFcY5ksOJpfehuiFbM/hPN/ADE+uTgEu0g5Z1f1cYN5h5cIdWV1+bQ5F
0LRGCqyzkV/jSlJAPU6nNr+gts+mkS/Sy8QRe3nXd5XniIEcVQ2nLXMS2yOfrgWqWNWQOmpHl4UQ
9k5MZVXmah/LnjTP/1o1tVJnub0sAbwECW9TQfDRLA2AYrzhQhsRpLncU8BAlpg29RqX6HW9q3De
YcBwwWCpPS2l2Brj9LHstfphgF7vEUNyVOWQSZPs/DAHqlssbLTNDObHzWTC2p4DBN4ueDkkhubD
t1Mu+BG0kBQ1hdhZ9SkJb/iGDLDNEyafbnpPXCYjs5ReUplwZiPlHTXGcPKnREAf8TKaazIr+TWL
GryTcHEuVmKNaLwD1r9syTsQ5ASClIVyxkSN9KVitiIdd7+Q2ZzGs3TbsXhzRQxg1l5aUmJn2de1
+K+aiaUH5+P3ut0uS+juo+m/Fe7MM0uaoYsKUamNICDg8fB/NDRwLF1GdOrkHDU3jr8udf90Clc6
+v6j4QFJ4qLi743fSOLUQV3N2FMYtxaueKHNb9Elx9O8yEflJg89c5riOweCiug9/TpU6GI27Udq
W5yeVuRSZQsxWg3P4Y3JKX1rJomUqF/A4yX4JajAaDxLfIIrll7T04k7Vmx7nh6LZbQIJJH+Uqud
qwFlJC427fulH0MwvARaKf4zZY6aXqwAJnzMrKIIIf0sVEM1CyWPt1/a+EVgruUbPAbiDyQOb+7V
vkm86uT5srRc0aas5A5y1zhsFX+ttaSZhiq13stXIa1ktHynkfapnOGIeU2YSqoA/0fHNqGy7orm
clXo3wgdpgjqjL6LAVjqPrE038nfuC4uDRwzDe60Mk4IKaVdxlQKwi2lO+JAIJpfWK0Vvdd8RVlR
kRg4erEvQyT6E+O3ipuOJAfuN7hB0ZvvIcguXR9QJS4OcHStyAE8gGO+Q1W650fcmZxID1k6I01f
T/85m4SX7Pd8+bibbsL0cqRh51YmGT69B/GV0dwgGJ5IIWrbs+ab3Ae9GdYU39ZWusynqOMulIdX
ozajk9psrxC/G5PWfYkAVJKL1AhIMWcyjVZN6anLOUVok1/XrgKBxTDkSgH4K3p5pLiqeqMcsDbR
Pzuu0wA+6PELB2NX0Xt0K3N5U6nwdyLfH57mCH+N/H1Ys1lRIo/+uEEAaWZij2dDG6dtherVhBwK
35qDwpgMTx+jpkVV3+jZcji1llnGTMp66uqT/qqc/O9Zb6VLuCVX5286XL1FtapNNA3QaF/H/nQW
r9riW7WuTQLOdkI7+e1MlyoQLu6uEnVQY4xhn8nK6sXvDGOLTesxbxyGmpY4q5yQTvHNkQ1uWJBZ
j07fJB6/EF9lyU7J7WezECoBobJKISlWd0ZPKvpHDviXIsMfkuqwnUKp2YzKBk/MDIiAHfDjNcZL
nLRbAutQgJ2edrYNjKI49fDdtlYGY++WR29mA7dZ3U27Zvl/F3RlT0/S6Vvhncgwxb3iroKkHVYu
YZBtBJnKjLPrC6WIavlCg3Na23YWDpfCR8vOq+Mr7A5pny0AWwqB7S6MNW4av/0ZhEAHJdI8tGJg
jdrYP+34gqJYyRZnW2V+vz2bkj/hV6Du2efZ9av6xylmu/Dq0PQ1AdoNpjo51SAOEjuqmyMbSyE2
3t/9+vID4Nbama9Es7mEK5MFgJo3U3aqfTW41xzUWN7Uzvqi+AyRQZsjkg3nkn6vCzgIRZUiqzJ2
OGwZSVWDqdyRmWpxiSATWeprkirNhaTOy4y4xdymeh40afXI0LqalFY1bHqu3LRIoQNMmPi72OZ5
xRTwZJpwoJ5y4uek4oJzdYTWrTyDkfYDMIA7fT0Nv6FywFeqeFPAE7yqxzWzYjUGqAYLLdPTi6Sz
S3RMlGcA3P/mt1rcM4EfA5p+6aQs5/NjW9nwUjyamLZz8bxwaikb7Um+ZyFHlsqU3TW0W3Vx/6To
8gr7pDWCd3XFNsruIyudUTikgSqW3TzlUuTfhOKlIpQL680r6gDiLy4jMW26vd8EtGNkEhJ5BlI8
pxVCbhW6KVtHmFgN2o+uvnOMMdZB0HcJlRAt4o7mcp+r5WnUNeA3xINy0pYFfWF86ntr8cNHe2KY
y0M88h3KsdungHsKOu3jbPo6UceAkrY9SF2QPDn+Scn0uO5PIvLtwYzYkok324gcViQaynmO23/I
dksqGQJlwh+5rdNWknmWWoBiPzQ4u8L46/yIyXnoFRMRbwl1+jOpEor/vuf1Fkpx+VRc8BgJC6mQ
Fg3iLf+1qUpRZOibZG8OrYnn0EoXV39ZVQ8Ke0IVDCBFxtMsCfhT9655pvFx21kq/9nnZpuQRZx4
7w9Npq0QY/4cFrdGGkiXNMFK1RJ07CXYgJc8VQk0ucQYi8Pouk8rL1hg5/8IPewxhR/wiBgy2pWN
Ou/Ove6lXl6SVSA3Mff/xP9SbfKZTcWgAaUkXx2Lcj9bOnYEMNwtNilX9n3412+pU2nGeb95CwGp
Ey39T9nFxXGZE3IUar5aRZYYRdVNzsu9im5tWeV3PqsUdi7QzspyU4eyB5/9K0oTNK8q7sV0XNZi
I3jJC1rlyWLD06DSi6mTVPNGWlyDdBdArHD1K6cVsh4gVc9/M1e3JLYjULbiDPHXaozw/agCpcyd
PAF9RpiUEV0K2vzWF+kEu8fvIi1zHDx5m+Pg1zuOdum1bniedW+hyb87YcRSAX0vPABs6Kw26Vps
MDYn+9bp28QGnzwzyzWIikJ3yWL5rnZ8zQM8jZ1AEIk5s0qcq6w1jHkzAHWEo7j4aSqZnOzHmQhk
SxUtqI+8vQ5PMPCX6cvOWiv3Scc7hOvGqVUydqs/7TXNbe9loOz1UcUtO+IsXTgVlmOwEb6K123x
Ni3ZS4clpHS/3Y7VnYpWcU4g5ADghKjI3GkjS1rpus9HAYSqj9Jm91/s+L+m3lVSNmCa4AaL/Dc2
52E83xbMF0Gr/ZhqF0U9jbwznWk7KsOoFBbqh6RWPV6MEKj4ByV+SGXd7wMeRkVypOZWmGCKEgTM
8k1dMjiCEyGWx8oCQ5ZI/Uw/h9QBdlz6QbNS3VV57CQljZKg2dVz1H9DsiO9+jQyKo+2tysFpBHo
f8P3yxhBCFkAZ3fw+moiG6G/DgVDp8alTUjjCGRY2XI1/NarAEsV5u+NZfCB0tXsQev8NYLSFLNM
Cj4Vsnd6hFm7wsoGDLfZyjAb6lyO8hVmbXu/2XOOOaKc6jcXN8YSni10DQzgNkD1RN6erjFYcgjh
bDjOQ81EWZPfi1feiu/knliBYwRbQ4Bk/UZfMWAOtjnT5K2zeBgpy+2bY+SUDSCMROwkOsOvg0tl
5bULMwPi38gY4pGm1ugvx5befhiX8oY23XIhzgxE5ecWaRG6EzyKlfQurfibeGoF9zRwrtvD1jEt
chqAkFDrESiUudEDfa+ikVT6MMeVXBjdygBPqgJjGdJAXOJzP5aCYePplKDaR+XDRv4VcWYRHb4H
dt6IaFAaSRfLO1wdAXgwLSrR5KxSkq6Lwo6qRDwIvEgX6zjqJM5lgxbmUvCwmrl/a0ubp0NIA3mR
3KtA+aN6SAmCOKyKgHP/KXwozdPWZ2f67/hM5nU2j14/v+eSsrgSTaVZx/Byb+pMqLMNvn19hx8f
boHIB7Hf5DhqlZQXo1194P+X8HC9PZzDgawv+x41ApEBAIKnFeKMCgOuDgQCopiN5soEim+h6P+Q
7VQRUFdCqEMMELEBiD7b3zGw9vHGxsrVYh67KOPNWGZfEqFEKyvDTH14CMcsMvzPDi+jgx5zCqeA
6VJg150Wn3Wn8QOG2bJ1MBEVj7Xh0xYBhP32N7WE5F6b8Tmodcs610HpJIVf8rJMVPSRLtBmHXkw
CAj/fK6qhcrBdneOWTApFzJMCpf1/SPQFUac+viiOwZfLFONdZZaGUNvg9rHRpgx9FsqP32OfC11
H/EgyndfqkrqNHCcQWlrNSmkM7eqAF4KWOrCSC0fzvQqfTyhE25EAEtg/hhcK0+C/BBlC8TlYrDE
9KNLjG35B09+BIr+QZJDb6e7RSP17BbQD/S/2H713vO8qYbrotjQ2dDtQjyQ67/TopG9VevPYI90
IvMc1YmYHQjj87DIyK5gpuFwv243fjktNKxf7TFjJH7LLXuxRf6WgVTuS++s9D3KltVv9x8cZCQr
MqsctwF5n0R5gdGpHvssNKMLbao5TzAIpFvp4xq2D6GhOmz6u0R+/AX0qVIk/kv4N496VazR6UfG
uvZ3+LBgUo46pQ4q5orywyGnWIFv/sGeGjcYoY3gxnHdLbUYj9FVadtZKXQe7FfMw/+6oBtpE95d
lSc5GSFFwGxmG+fKm335j7+u+ARE3Eq8Mcvizb5XPdohwTePPGJKakc6Dt7cif2M6MJd9mdgxQAu
kvr2RSfqEughR5WPFAe1ouaeUSVhTcY8VSHgDn9ezp1692uODsSOu634HDU5NVmd9Sp7C5yXcMJk
93jEK47QntZHLNl47rct0jq5FQuTynR4RtRuZjK4nA2kilSWJfbFS5U3Y6LkCiJ6MHo+e4o6hult
EYAunPP6d/124SqwSqt1bUwTKbZFFS0pMzYmpcTohZ2Qc5MK3muPOzOmRhuY9SCza8gYchBPI6pe
MSVvrz6RwUaGv+SjnGXpfby4fRuv0FrjF9Y2N7WSURlXzJx0pNHEoh0sd8QLtRd9X8JEVoHnHyE2
FXiqepDCf+Ziqq3/3tClGjEIzG/XL6Fg/UnHMgAlY9DOi4KXFnWZw1KD+jBunIDbgzHlZ2LpY+JU
6IPdAiskZR4WcQXesBvMVKJMeuqh06AyETOzuQqOyw62VZBNcWbXczxjqy6o6OJaW6rfcLcsVS3o
prQpzPNGk33RXAJDrTfbrpnQtYY8pfpP1+cs0PbinxcIFRi8EubZFLdmPJYTjUYNoZ8Hu0jnUlwX
35DOpW5Q33gqg0C2GmtU/vIzWY70R5jGTpqNPAHpzUCpEWRPed8FbfhSQ+WvLyb/YX3uYH9SeIq3
A+DZ0WsTAZqjPhcsHH6DzKqH+8czXefGPtCswZ1BDtGOUsbQ1CF636GSFnYDh0S2iRkgpqerjb5B
EK3sJp+tjPkyqVpKGx9/cDBkZU1/QzC8JRHYQABkxQsFfZ/yP36XzaeVkcju4A4NorbE9HL+ihJY
RmD5kB2KABfycm+B0w8AhFmrWi1R5HVHuJWHLQyk7SV0FbA3UrbuN0W/od2VpGX63Y7Mxdzdjd/+
j2Ncuc+06r3tBDNqf1+5522nVAecmYZDzH9Qf0JuvqukzWiP4iQMjs4aTEnQuZFYny+Wt/4hEvor
z4maS9/8NnBFS8NkmwKOia4qkpY/AZcucySkB/qNurjoX7cu1715+WhV79AQIexFcu1rM89FoEE4
Uo1hnN6rHw6d0tyU5+b+2NCzwpU12sNhtmKurkfkaL8QxHyVIbqf0j6yJBFup1/jHS4cRtmvaADy
3Jv4+Ek5gMT0WGRPKNY/ZWp3SPOSv5wuZNbfrbeoFh8yGPkX5NJcsPflHoZssykCI+C9+68/Z9cr
lW2kXYVt3wJiAwr2mL13alRJdie2NUQOxoP29chLk1huOixxrV3AP+EBZ3w+p5ZhHH0IbcUcn4yQ
jcxPZXtK6SP2g3qSpmOHxzBVyMm7o64OVOMZpTH4NC8x1VvXPTFP9Tlmq1DoShQLLTq3Yiu/KZIg
PNMXg1dEXkiVI+OS9IH5GIKuOjgekTBbJzRGYk/gsXh0YGkx6BDBuNKKp5FUfUx1jYz047vP+P6u
deM3QoHzDs6VcDSibHBm2An5hIZsdNDo4y71OiFqKNz3xGXlJXwkxd1xRK81Pv22reqMkPkGKyfZ
O+QHmwUej8FW2GiXywSAr5j+JyWz1tBWe9FxTJZ17POSdm2Y6n/qVmFWSl8BcnV9HNp8NrKiw45A
xtipwi0dixr3TF4FGqB9jB64oOA9b/GYWs4tJBgqEbcVw14yysZNy4ft/TTCqJXEDdiNxEYVIq8B
306E5S8HX17U6BAQ81fx+Hrd+656rcy5vOm16fm+XZubn+VjZAK0cHW9qc+LS0tGyxkeyd9xMRG5
PbOqIVAfghYSTqDgdfU/4NQEBa1WwI6tSoy4LBvn3VX2+B+sd/UbJWlEeHz2NK32pqaHV78W+WDo
MiMEeAIxEfGWhyExvBGsCcpLjDRf3wTKW586f5dcT9ySW4LEXKm9VwGcE+TOc6W4f8F5jf0PwAR6
mR5mNIQM9ONJdW1LyVVVVExzrYLpcKlTYnKcq+tEK/RnxpjiZN8XPFSSU2hVP+sjpEKe0axX6sjk
6F3OtveXZPuvh7LuoqH6QlWQ2OpR7mtEIQ0LQdooT16R1n5FfpYvss9UOlii4y2dDdTvT1BGtISn
9UlNEqkHt+0TyWOoZ+BEsXBiSccgMQrPZqbg14VlAvsNq7hUi2zfOohozAtsDxDawuLDOqSfFCL8
VEBvEfOl380ms7x81DJ58PaBTv+ftHDbi8FU8pMBEVS9Csqx1id50yORIY9eq2XHUeoH+LOuGHvZ
7g+0qby434sbGUb8luXvEFzM7CJobN2tPZgUCrnBV8xtPmjMlq3Oi64Cwe2A+brwYe9vO3Qs3PUE
sHFafuQQcUJzAUjA9g5EEiK+P/8LyQF/UpLqwgJaFyQ4heqfe/WXqNcrydXG+XGNgoBivmD3nKEX
/DQsh9OtuUxRIpM71XzimaF4UsJqujbQRXHBCYn8DSwoIBi00bnKiwy9bD0fq+bJrIEAdjOpCGi+
XO5eO/1g6/I4Mo+xcd903m7X34DdtSd7uBp2Fsgz5BDRKw8aRTzj0/LfLwMhGssDh7AfCXTIOs7L
8Xp8+MQG1aI/xTSoNnMmWvscYJl+M8YZGFv49UHwxakjlkNGgBZhSBZ77KWcvAS6YK4hwtJ/ejSv
ACo31j5Dvb+tM+UFMMBRmoy/g/eemq+L0koHarrAqLp8Yk+TdT7Fdu7gC9v7DZJbh9RbdbEhM+AG
KvIzLtNq+BJhKHm7SMpnlIsumuNC1U/eBV/R0BY9jsUqomsGrhWb/WmKGQSI2xUCA49yFdfL264i
3dXjEIbbjJu2ZqSjF3I2MeNOU4QeQktetZC+oj8A/15nvIQa0We2+1VdHAIhwOsxbsNVzuhdW1qE
c2U2MJFNMyQqMIfx+6PnlZRT4klt534zCKZW2o/nnHmiGOhI3qAQ22sF0q5S7kWlm0frYhMLEEhX
MXnl8mgCQLRtQXsAdRQqhk4evXuosF3unzLJAHmV8UPx7peIT6Meiv1jKHE/Fv1LbvfUpUaO1P2V
Lhi6TsIzl2LV30e9x6oaxxTNVAURp5kY2OZD01UuvwyvR5leHQi5A3Jx3iEb4BtOcKx1019xI6y1
NjuDh5N0ae+0jKDayCdZAZ7B3bIInlnobiS0NHPkp0HH8CPFPhf1caURpUmnjL2CdlScSxH/jftZ
61ae2WHozVuEZFE/qz87hJT0y3LAnA6SmJKuJS9mW74v2nm/1+d71YgQKvXl9KgJqa9gZLXJiIBw
at6o/hyyFQXGb+sqmIEYrjJnoPKycpcS6bR8AwY+ET4Go5XmmhKeeylLhuTHOFY6MMj1+YbVjP7m
yEelFWNy8OQfMDSKXebD1/IpCDz0HITa4xbdiWWy+W0aRdYuP+zXl2iN6yvlFw0GnOP3fkx379dI
kd04w+hHHiU+VTZrwUfk4opcbBNwVX2BM6YTQG0Vv+njgQtBMo3QrFNeLV55U9szxRMkdMeAxPQE
lQo6RIN431AwqGpK4BI4+BKVj3xer2AtAyPB3RCvtbNjn+R7ldZwWlZ3pAUaBDwIEdZpWarLMkkP
65pvx+oWpGvHgb+UJG9UaBjzb0PMG3spo/yeIgCcVFE2vNXDN/aHF26eFxWEZKg8j/53pBBFnCFF
b66gcZslcaKgNubXLRuNv+Bms9vLZT7zAoCgEHa8FGez4PhA/ENmwKuhvo57kNStGMWWVZLhckFq
eBG5ByvBR312OHp0NnRLcn/ZNmc46XLVzuqc/ByE8b3Y4Qfk6W2t5qKSKv2VBg9/o4v6gpr6NzBb
wsc6EDo6k7g/HtUn96ta7kUktWAKg8ZgiiRldqLv3eY75dJ9+358b2NvxT252wyD6b+5xFJD4LLB
+RUm5QGEy4LYaICP7BASG+4rg730Rgs3b611DT1YsxgXPaEWinuvXSb1ADIijmdWTZV1IACAw8pq
tu17tuCFBiKuqQ6nDDy6ThV/U21ntrYau9Eniln8ppd9tScDbVEgiOQYkPRqvx9vW2X24ZpPtGpT
hNTEqOgxgh8qXDR9V+ufD0UUKQEQN1MeEbv5u6SbxfR6UMh59yi4sxelJ2ZH+YMNhz9GCVJRVxD0
iqyN/8jpvhCChMrSQe1/7RwfDxOxBERkfenXvf9SWoRpmbWBo0XAlZw/inlw97EWmvy8LUcmqh8K
qcpUAskHYEHqc2HuEzc3ZRaToeQYiE0q1m6Gzt0pdA/17Dtptb4F68FLBp9pvj5pifAmk9nmDJ48
633grKdUX1MFYcigWpcZFQSJ+1Po8odhZf19wWN+WdvQIL0lF8kT56E3AelxoihqgZx+p59HjLTD
lb1WEZ2esQ3feSlixkNyFp7fdumbf0ay/uQf59HFZ5uRaOPYqfuMrPLyGHoNUjg7vFD99LdPww7E
IxBtvDvzRmDnEzy0kQW4z1vjAVg/FmLz/6PgICidYLFZMuT62aM51DGvmV2DLwJ6TMGh768triN7
WmeznbkDQyuN2Zat6RHWxrK/UYfG0LtrzcG5Nrw4StGpIowDsAED0h+KOXNemP14B3X5adVPZbmZ
9W8bNGRPA9g9fyegtsSCFnkvcuw9Ms287ZzWoeQuE4Lutf8u0+bBe+h3PCP8ltu7hDAvKcJqdREH
NA5qjYPWm4ru2i7DeGP27aPGZxxqPrzgA86UYG2YxJnPtXrEvO1g1afKl1F0f6AUppwoL8lBDkPd
s7VwQCqVNWuiN6bLhHHANI/EncYw21tkwbrHrlHvG6jm/B7mMVwH11rqbVMWFnwX0hiKcMhCPb/A
qksSB/KXhjG6aC3xEiJ40ysbgRRldwKWVOSK0OqzpeICntZQmFLEjJtvwkm1jDQkHPHx1fC7P0HG
TutN9hRBkJvE2AylPE1WNfhKMBmCnG1ltMl8prJbHzNqaOLfBc0yBKZw9vBmhujXULE3qtiMEJjl
g4CyluAZ2eW6WJVvXC2sK8qMd4vsUH0WYsWn99KeNRtmR+qX5IC6CBSzpyTgS4jO9wC+2qdeCWXO
+SQgQDKzEcqFUMoiexQxVuCvB95hKvgnOIpw4uprm7Q1UdAxoDT2KdDwJ5uePBeW3a1tV2tmUhPM
gUR/9FNx7W9Cu602F3I3MdWS3d/J69XnOilqnDIcPom1EKkCYn7TIRRg+orInBpt/FHO70lNfTDz
JsO4/8CkIC+dPmUWCJr02GwsnfapK4hHSXdEF/2rGm41Xu/Vf6QNXqAnBKHJFnPOvrA31CtGD5x8
f5X/5C3c4mUfeMX2PwgAr5K+EqX5ZH01yj21D0pgoId2KT2xhjwRKrT+nG49VGCMrvKh9nTiipTW
nnydINYcruxrQd9e7k02zx6A9ldltWLKnyqzfD0Ysh+v6gpvlFDK8Yg54+5eoYGQ4u42QlplRHxt
dBeXVuCSLqtVN3P5G7W5enmtfnS6iptK/0Vda/ZERLc7wxjM2mfBtvvUvLphDA4W1vF6xSq4h5Gd
7Ib+frco+ta4HSIR/H2yTcHSNMzL3cuIEDZlTjOhhcakMoQy5qNXjrqYboe0eczBg8LdX8NivyNR
L2la0a1OfNz/xCEOCFMF1U+kwfY2kTTWBQhthBLMMrKlcCBxDAUcn0Pj0cqByjsDO9OKSPNPHGTe
XGkz/0L4Mthp/0vyEfpTN7jk6DyFaK4SN+B8UIdP3N7+ewho6QOzES4Z2LHEQ3LevayJ6pty/y/h
iOUzfmvRNsf/Ozl37HpeAxrxNgicDiKdRB/z5hQKT6QG6TQNEGMnPBd7/rTS8V61+nZ9R3FjYoDs
4dreTqkllTusvnjSwBtyfGIgB3Qi6U3ORxWtYYlvyu9ectdcfjSUInfIYMZgfTTJ3sVkNw3b23r7
XN+zb+D3eUWZPaODJGuZnGhLDpb7pJlYok7BRBkDT6XhZQ4iNRbMUUtRbxvMLXWGQbN8Rabhsfx4
FfnFxy2kZml1KCeJ0PZf6cfzRQsYSaNqmVJgX+PoZ+2vlJIIN4dZMTXp3G4PSus3l38oB1ruOxHf
wOUFlpljly0BpGpM3Uwb/m/+tOVctUAwX3Y5XvIz0HLc/RJcXY3RWl/tpynMIi9hI24I7WBVhHQa
Qy+4ear8HUiOdtzV46EGDSQ2J2hccJIoWyXS7jC+pmkxmSzBjhhydmZiMdLlqbRKKbpgUlcuX2CM
hfkvbPDLjwq3GFeordy6O8jorj9lbvJrcZnQuGWpfCksi7fxRj0rp2yE28JPnanOvNNAKqqUm1Tm
XX5pERkr7RNabrWzuHV/fkxK/W66Ezx4McQ1SrLGLOpYSR5y0QWC23WBoWlt8pqvYaGE90SUOsbc
kMAZr8jjTAQBN0LI9Vtmv0bb2sHIamYKVVhbx8wIwvA+IODwwqO3aONj7S10KhDr08UbE6FJY77C
plfOzZH6kWTZtxKPDvy3A1LDYdWi9ZmrwdEKf/z/4+2+uraZQBC9tZl0JH5xJIIQER1bBdxnH3o2
jSNOigfUcqAZedfqf4aqWYEe86qxk/b1lI7lnHk/ISe1S+jb69FfEDBYSGPQgyKiuHp4+oO6Qu8o
tu7zxfE6uN/2NqlfL5QszogRc/76ehdqDpPOyj9CWcbfaw8J9hm7FiHAv2S6koroKkG3zZv5imyN
Bs/iSUz3cGr8JoUvOBuQ8isVSL+m3RBiMm+/Fw+nFY88N9lYAvYFo50k5yliuj64bgLCiMb7AMXQ
F/3vtznPH7lKp1CQa8RVUBtOO3ElN2N7GXhspG0970VY9K1CAh6jDPgcZpbQXzCkUYbXQLr1uN9T
HBFLcmYHGJ7FYK95V061+Zh/jCpwBEYhwwAxrUmEECXpCVhSuFIYbkFtEfP+dYN7ew8jCH2Yi332
7TRGF3QNRgRWsAFdDes6eVJPVzCd/mCfd59jWvwgL6cqTur/mFSoangx/RfbfZOmvXHghZ6JoEXq
gOX0Kr1qjF09vJBgSsj49M9rqZcHsagWRTDjlsJ55DwmWzAREbU4oEIEs8TjQezAWpHQ2/d+u+05
VymrTk3zF77KqM9ww8JkGM+iUWy4d1dcWWfg9SQd7lCRkfQhIGOfPEzE0PpqxSZm6/xc33q2ecne
eOHm6jJSrSjJrprQuexmrlFRI8XiQ8ac47zB7Fdl3ZNgHrBckRhNmIKNJSPn1cnxiIAgHjj6PyF6
AiNguzyJOgEbgIcoa1oMMlv7CuL34g9ZcMEDki7sNWvRZY8HVZ3nawOA+OqsZTArd8Gn3vjDVm2k
Rfl6Xbb1OZtdojRc/nxguWwC/TKZYbAcS9FgzEjkYs2FFUoMpoEhwmKJPaDwog+BbBIF+Qkghbtx
CvSZrrbGk3tK+pVOXSN6sDuh+53guuPGzpOUkm3MUm3Lm6/eErxT+QPGupBsQziiXHGiY2vMecf0
/UO3a7w6ePFTS9FBdugn84fwQ6UgLzcXD9OmXEZM4vfLO21vEASomKa6s4ZM1wDzrkttzDQL+SNR
FTuDYn5zhrKFbU98zQpAjEs6fFioeYu+On+uonzOc5af4Qyow78JnHGN9IphoT6z6wxRyeBiv0aE
p7+cIJi5bF55+V4MvNvmtYHU5RlpieMeh8du5jwyD8g9dahvxtqlHhugq6koBumYWQYQrkMSoWiu
w9vrLCeAHAcppw1pm5avMGTtMZ8zlb9blkpiGbzG2xQqFXdC6A8ZnQyMoqTrPjE26OaQEWnF7/Ur
NjhZXPoicGLrhxo+G7/CR/CNlDeLK9HmWWHQcPh81oLtfouQtZAkRTSDt9jOlWzM4wVS4s8bGaxd
X+5e1WlXXRO/5Kc4dNL7W4VBFl/hPR1THRe3chx2TI1qzzfSEegGhFw6yCBiIuvTQORhUHqgzZqR
hwi2ekj7XYcOz8yUxmQQObbeRvPMPAIKb+u0kg+8RsVjGMWBYkhYvGh1g7mvCTXvJ+ereEgSc/Bk
8lw37zuLRJ3Yzm/o4Nv+WPN8x7vL3klye/vgfAC53pammm4R0EYIRgcdo6OuUGwC72WUd8T5qfFS
YYvWFx1JKOsZaV/T45ZhMIyNuoGq71EzyL9BbP+nzYIzdyHUSRk3y2usgHI9npXZKmK5/mZ0xeYD
T+7WWxFtIGpKp8eh+wsWbRxXatzxBAgszUjRAYz8YEhhyB3z496HGF9xajbh2exU4lPjWdzNvJr2
JibH+jLUxGHYARzlhV8BDlidiQGaGe6m35XnJrFhipai2mmh5ATBVvbJrDPUkjXaCyfs51Wxr9S5
tNJZz3edCsU6OuDhOW72YVbA2DWtJq9QgF/DJVPj0dPFQbXD5fHg67xtztpZXuuSy0aRhcQXmoPC
1D3Ay9J2Uki7imDTHriFo4P8j8xukqopNLCB2pzYZc+ZCbF3gte8BN+zJrAppdoVaQNdYjgi3Q1l
mNIcmxI4s+GDqRbOwkYBDcbcnWeOHgHlndRY04eQNMjQQIZf1x6VrqHl5QHWrdtcjtL4b+964Dfv
FK+yzU985wQIcmrkynZEkLntZ3AUEMuwRTVHPzixm8jeifAYG66HvmMFwSrkWb34/UnR1WxAtUw6
yN0AptwqeqHVmhIq9GwJmyou434179QQct9ISEaLdhnkBTpsS0xGrclRSLM6c3Cw7HnF9kQRryaS
d4tJd76JkYmOoeRh7U9tg5jKhKsZ1wioUJkvURfk0MRQe1WqfWuHgLx6imm3qUDrEN9ZGl4jO/lJ
rDIOoMxhqVFjF+Zmfmf4MtckM9zDKBAzYVAFgsvqdX2lgeAOAfxzTcqtMQoCP/5mqsGzya8kh4Tx
uJByJwG15tn0csA/AIonYmyb2Kq/HuCdxKyDwffJ5CgnTEBeCmZGP9ItVBdBaGuAnifhCQKwyO1i
GZJbUeB22OVueGFiSFb5Xzm42ayN9uW7jIe36qiWF/ADCE6GN5yRnV7iqrZOqgS3igR8u7JkIE1i
PTiQ7R0Mx0F8516HA5ndX7m+6rCMu9Ot4qMuvRQ0XTBP0mA3XlE1sv29T+hDchx781rEE2pFecly
m+haV/7k14o2zvpqHjVqAiDACt73ZR4yVW3qrgfg75MaWpWo3Sn+wsHdZJileHTSwjyXD2UZJlMm
ZnFnPQF+OLEZLPxH4xUS9PXrECv4Vc4M2oS12mEldNzaAFpx20yNDvi5TYNd8n0U57bGmdd8uJU9
Wto2sD9F8XVV9rxG9b1KT6vbTnYRMbeimPVjggkLYVubdL3ZUIXP41XQ0aup9DitlWFoxeYibSCM
iLifj0HAFrPElvBvdq7YaLLvN44XCiqDkBqQUez9CvKbsGuRffno8nVb+k+bL1Sy9+yKkW+KNytk
PVgBq2g1RIhiuzUzmPZWwpKS+isDtMCO2ESytOrXTALpIWGPrcpFpzZmO1s2B2Uc9FonWpdj6u9R
Usf6MrZRIMmejbSDYOAYIGkFH5fEg/QXULsZP9nAe5IRN/9NvKEXWAVWgyKSuIh0a452BW2PwE1w
wU9ajFfEAGOVSv5oxCNqgy+aI04CHpfaO8F/stumKa2M0GrBXeABYKFHAd2vlAbIzJ2BGOrYs9qJ
FqYIWRVJvDbBfTmb8c1ghI1XfquW1FSeaYYyNDjkkGLW7IAx6bg6PKTl4TGCjbHXRtpsdJqU8CHS
A5ltG+zPy2ev6EVL8nj6Avet/SYSh41MYgoJuyDm2lMGgT08fKF6Bv+iJx7XY8m95KacqIlrAIkA
Z2KWVWyCLJpIT5iEfO4Jrs9veaOibK0Gg5ZWwsbNvPLVYAY+c0UBW5iIceBsIVMPupd0abprr3n6
fvtPs1+lvIAC0QjcE3hrD2w/0cwiuFKOGMpze3Xlcobax3L6/l9gqBTVEGSPvIokQXyWS5YT+do5
IeFkUykzW4SCAbL/3Wodrb+VvLSk8Jrm9f15OGXAtjTLENL3ji7e5biCF2T8WNIEcDcMeWmDBZ+V
cDC2+cS/G9V8AK+SdlHEyWDjfusWmzIrZTpLR8eQ5ZHXBHlejVd9/MinZUAfoaWhQ+CccV2MohTZ
pTdRC5k8SAYI+sFxU5FXIryMuy0GW3xUICA8T5xoMuB22jJekIyI6nIzJfxhn7IIyG5o5G6yWVA9
q8yV+IkoqmMkpMLGW1LJkYL2w5YgM21Iy8QrJHylvDCJ8N2ktBZJQwMR6TDY6RrhbQ+/zBGSbZjX
Hhg+TBEUeZQF64qs3lWeRG4KTdoBewXjLFTHEYQ9GZkxLPV2Lr4MDN5fFOJql45K2hjRkI+Njx8n
i7iU/j7PQlLLxNfqa11uCm6A1FsNlzHGWeLCKxPBfXd5xuM4o5C9HJrCMKv4qQZVnSUPHFYTLc4U
15PeOkl2Y6YY1U3kWdKjdUHo0lhKFgpzDbqnfj8LHo3D6QIrGBKcB+OKuM3399N4pd87oE6u1sqA
8kbNbUkA6C/XAlFTYW58eWbQ0yfQ/BGPaAees8Yc48jRl4kzlPbVp6EAXu/gqGEJaOyzy7bKMPt2
2DQBWIdAJl+le712dwIWVZdgPxJyg7jB2sCzItlACd4X0Xhd2hQnMn2OmStos9siNsV8XbROstTl
v5EN5kk3wl5utgKj8D41U611tR/Pp+hXumwn8hc/r/ygFX/hF055Ks2+UeS9wyT0nmqVHefF7Pt9
OJNtqBWt9Vv8K8My0JyNSOQ05P6/hAUY93ZE1Js10cVzrP1GrsUsdzNdgJpyeuE5elvDbv2B+PY6
RIWW7MipFNxh1CBEFPcogxrilvAkCtRU4yKwqAuNYkrqO4PrSBWwntPVorFmDDkW+ZXxz6AF7FBy
oJTsiunh0TrT2IEFf4vx4wW3ZeAUjP8BS3aMCccGAFK/qaWedIJ+T3l81qi6Cl9HpaPFhczawmNK
QG/jkiTZwUoi9RVtWQCgDcbewtN1wAlb5VHUlet9M29BUn2I+2uyzVbLbZJ01oizLSCa//rddGkT
v4d38cuO0SV4kdIXjsaIcR+CJ6JOvLalF4XW7xWhq7eZhl/bLQ048USSmuiHdzH/QjLOwNed3kgV
hLjEypoxEtwODpEX5VxTQ/bCpYApqNIoWAJJtXP6G2mXe2MHnBOOzF+C+cIWTkg1aq7iy+L3R/7T
0FrwIGClH8wM9ajtXoF/Mkx2No+0AotsWo5wbz+RE4jIEu2gtJ0rgYV16AlW/ebiv8VgrteWn96U
ybRNLeGzmoWLNGqQtxD0RUkcpGnnv9X/J74BoNeGtm0ZtvmbsmsPeExP5CudQSp369/q1HkkImwj
SPJswxFpXBCZ5jObqA22m+vn9Tx/2H5hgRDwQ2bNAeXK5bT/ZHhBhdqyGRjSM1rqlZBadaCA8UiU
SIyjgVvUzlC3u6Y1ivOX6jVc7XJnD+Uz/EM92t8SG+uXdCEUuQeC5rB9DfEROPEmXcv/r1r5p04A
bGgIbZG3LLXgiE9VDu6JCqwTCOKe3BTmiBMiezXgR7zPuPf0lyrakkKCaTOml4wfQRaXQaVbZddr
qoQR554mR4CoDO/LugZDlIfz/UD4xRoGwLJYuRf+9flW1BtPOnAudQ29KMup5fBBCER3Fy6ldTtW
sGeKVCqnzmNCc1N5EPEz/kaSxFfa/YXvKQhSDJd5I5fjnx3uD5YDvdeZaqW7oHEO14L5zHdJKkon
shE1FPjDYSmcGPZ25tInB9uqXY28Wphm1OMBFWCFgEAZA7tudYFamlBF/CLSzsLr13xxMH078g/2
ifepe22dH3edxn39onkFksmYQ/R98I87+H/5V1BTW8PoPy6pROnW7ATGvZ2Fczw5xm2srw344/cm
QuceaFj1waEYXBBH1LinMAUXnXh8CgX17bX8tl0RFXP+yrvyasO4wlFrHDx4fe8sCs23lhN56xLU
ohcD+rMz6J3eT+sKlXmnjRDtZ5ieq8aWfKN4seRCjDu8gEN/k2luXxUEWjg7WrHtyZ2h6nzHq0Jb
kv/4xDDXTbbNPTkZXINfFOqN5QIrT7oOn/272KmSZtFahklMkmsmqYeo98aB4Oy036rDPAkgli6+
vx/YVo7QO5dxOvODpWDO4Kv/oYgCZCpwIa5T/QahoUfIdAwT9tJ5Up+vugZ2yRufq7TpcEGwG9eO
i7OkN91fkIChR4BYmIITF+xdC7gnT3eu/xIGjhMlCksW0b+9nUodTIGF+qzJi2jZuxfE7nVaAhjr
4kQFZRmIZMT1wvUJB9hpKjaTIJWPR9AqYxhRaCoZFSm6C1wpykFXM1afX5CqKrfjQfuxhvJreWJn
jDxazTgLcC7F/XqrhKssl4LdJMTqNdnDBi7eKe09dcmItVTZVMvzAHFKBo7VXR5VGyjjpWNWP48y
gqYOHub73WxCzyqcHIjPI+VFkajis6Z78W7VZUAkd7IQU6ZoONLacoyu30tfnULif/U3UUtZvZ0w
xT4D5vUjjmYXGmw4u4hdp8xjRUFnef7rnhMkemiOV1O/ngeAxQxAbmDvCXC2llYyJW1l8CBUP2Tc
UG9+JnfTRGEc3kAbp1p4PvIVdzvzhLtPA2bhT6vjE9FtNHbdge7N1/2KenFcz5VCCNd7d8DIKnPt
hdF2aWd98QN6ycQoe4tA2nhkkYS/NagWjPGQYiehE5iJYb9JvoLKf+FCupkpgJJxQZv5lbgG3wRR
JfbWsqeiPWJl8+zczAdMPiD00hbdeeApBubAaJZfZeQZf92umBTtNzxyUtqaHod7wwBPtzztyCyH
FdQLU1rxDnP3aWnnETV/y2wJbtjKiS0SHlqtQjLO9dvzrPYfWShBD3XgisRIWlxAHJlCvUMS5Dwo
KPD1IwoZcQ4Uih7keut0/ecTVTZmfNv5d6lU3zUf73V5M8ZxOgQIiz7HRDIGOZxqS7c3AyFPxqhz
TSBQLiGKDF8nPC/g/vMnNFP/ezXYYuPNA3tieOEAPxrstfy6Vag0orsIDi38KeoL26T8AqsfK8M/
tmTFl1w9M77scwf78KxOzwCl/D56D7CJQjos+mlTGbOjnV/CzY0B0hBBtsMsfaTM2ZwaxBKdbfoT
oMqnK4NZ1/WmoscSgn4gGwGWySiFNv2eCzqqlKpAx5I4oiV0EfjrkuV0XDLiiApVby/GbUuUdZ8d
C9+78O/uDx404T40BfAFM4PhtWJnZ6SNw6Z/1Z3sb4MCXJTZcrmFMPXs5w38EVWP9SIIAMEtmvLY
JyVC21EId+ihD802CD4t62+9FGRppe0wRGO1AfrFEkeanR17ts2+7/Vvss/RTS1vQIaqcCtPqL5u
weDO5yJB9xf2OCK1TKumxqKb1r0nj1RNrkPGoVsI2zy6gprnB/NkS+eCBekM8vaxHz/Y+ubEbsZS
KkeFQrb7hOSBWqH6pXba3zqXUi8Z1Q4A3KSBJKI09LjE34lbTMKHZLijHkRIKPqHDtJfeTkJY3Mc
XYP6NFRLs8uIxnZyXpUEzx+C4YbkjLZM+TVa+uYrVOaIdf+76rxZRqt4YHE5roGxDMamAUx7LGsc
id9iMgs8uy3cthTyn6GgPffL+WHSqq+wqnKgujlpezhLelz8IK95Y9mgg3myjYj7W8v4UCqEu7kX
sL/Kp4LO/ooEubRfIPMwl8i9kIFbtvkAke+0iloh1SlHvfAj3A/BVB08Pi8x7ijCw/55l2a1s8a+
6XREgDkVK8J/Zk+YLRxs5AU0oK+8CJ2e8jH5rxe0uZ9EPf/97SmgurpGs22CSgds2Of9di8dyw5H
gNxr70ml6uhIE14CpLk1GiudU4JFVYWZ1g5/Kz8cxdCMLDHDjkOYdDe7XQRH1oGfiXX1BXi3WsrL
ct/9eezlR563TNuQw1nEUW9/Ei6x4z3fjGa77RrguJr2YTDAC7zUhBsGZ/PbC4OYpV1BQefcOBHy
y/q9crKfAkHGlYiJAm8NEfYxlv6J6CDcReSKRyyDKK5sYwDlvy5zLa7unVwVtWSKOhEzaNAKIjV9
fDWQSBtiBrOxP0rhQvkr7AOuFGA/slw0omyxgj3mDcvK/tYnxscE/raJ5+s8M9oUmpD5C/1XX/Gt
/beC2KG0tdox3INx9+QQhdVz4FaQZ+Iwav1h/x8/wnWFLG/g5y/jq+IJfYsTv49xI7BCjZfkP2FE
VtQg52G4RaShm3lwMOIT7o5T26cQJ2dTr5sYomWee5RKV3ks4m65MrDzUF/2zlz+i4p/+c3Hb15e
MxcCU2h4cJTadCPzwjC66Hd+XEu0C0DSY12AOUNnvr5yIXN9GdM4Dnqt+fLgOgKK1jMJv92z2rAu
NLYZ26Wf+05DCZnDhygRaVEstJosGsvs8zhskJ3DWLPiKXh83e6jxHVH5dq3MOJJRscEYhFh+zjb
U9VBTSZRb6cAf0aIbbB1DRq2SzgEeJ+JSKtC1iXQ3D5W6gPWgUAuvqALg0t258BeocbYRVZEPu1t
0+xqcsERkIssDlubyJeRV64aHhiJGg9R3BzOFwKBATVkDHif3YHvUcnPXzvm3fUPFekm74IxkC/7
cvGyB9BG7vQ7tfHCYbYnqKwCAYGpdcjdHX8NgXIgznyKzHAAuEJpsUb9LXLuHu+ivF0nikspsCnu
MrcXKZmHc3ZaqReOzOMLXViucMpJKZ9Kx9LPIOxAbPgu6lr/0O61LMaKd8dEiiLA6JXHQelcZTPL
xDHmSPg8d6M+LBFk4O7qHniCFl3nQOhowNZbUta56Rdyu947a6t6inZh1bZ0XR7YhvF9JyV/9Zsn
27rygwi9wTiNvZiRUWT0EUr6lMj7vsGMGyu4OLaNtG8+y0mYqeG7vxLkGGtK4+/T55JxanbLIz3D
SprFt+Uk7AINE7KCmqcC7k0DNULrI5m4g3QUfvm4ZOQcT/T5LGvjbP5Pl4xWBjHdL21o/Lv/AYDf
6kWNXpI2j7E1u/UDAFl1jNO5Hpu5KEBiKe0U/JHOxSoavCqNUr5pKyrTO0HWs7rn5X1hPRMJgFzt
pFjjpUyyQ5gbbq9Kvx5fZP74RpkDdWqPhAHynhQQCWFwPsZqSt08nRkGWBYFX3+SoOPqz7y33qRi
a+B+VkvRX9bUVuSy1JSfgy9aiigQJieg3IBtI8dSDixoTjAa0z17sCR4pOFkLhNW3Rnav6cZ2ISt
pa5ALbrehlt5Q+4Y0pXewAEdV2Fm4wc1NdEPWKkRsN2l+QEA26WCKsZFKl1H54F3gBD4HduFDD+/
24nphhAMe3h+FLjvinshyVq0fzUL7gvwlFy6fXc1zMKw0aF7OuME71K9UuTupHjlKsm8fBLnCz+z
TOS2Hr7j0wAx7i12ftCKOUp5YfaI8zObmyBdR11YdnJSKIXGYCbfDu/Rkaikut4syJzY5sSBElnB
6uYwwgwhTqtBJqO1y4FrAtJTzDnum37AQfeRIekCcfQFYIsCcjSaQNwLOl81dnoIp0Aeq9BWXWZV
uInaT5e6FzO5XYORV9uEcElN9y3OdmvsL90yHNQvnwL/dGHbCiBTdL4eDQEXh7lf+fwP0jpKrxHQ
FR/m1jclNdezWboewvixOEmgm964IeYR202FOYySv63GhzXmCPOV3C9dUJXkLJvhR9Usx4EXEsHz
2E4TqJs8uMSSsT1ZqXpnr93dIKlYj91xXA8FdCysa46R8t7jNg1nRpaXjncnsYEFiCJtQUxhu69x
pZjZbspxp1K0kCtoQ7iBMh9sXMct+ZDiTrErndyMR58kG0FSPu9rRsJv0vtakQugSllRo7ho+oQJ
pHEhxm2S2maKiNSSncQDxgh5Mr/NThyuFNe98QDnItE4C3dPM6+WqvetRtGoHGRRT73vlYYooiA9
d+y2uHBaoAn16Cl6k7TIqHA04MCck3y4Fj+x5KLvHl4kZ00LxtNQzTGvRP2CThbbNr9qMF/5bCy/
prv2mUv+/lGhHfrFhUDB51iQVUzjBU8UVpkllmlNWfOvH8vcNmHG8ziscb6ivicTeXziluxR9Jzj
5xHaRvVjpzMYJB6m+BRApfcaiStt7rwIt9yv9CvyZIFt10hndBoZ68u64AYXrRIRI64vdFI5gdYR
9y02d/x2SSSvsiO0g4naifKArrHQDqKdcha2t/o+l4C1ACI7g4IRJyRDD98WH/b110Ulvb/PXD0E
lQwA75tp3aZ7k582ZqnWMaOwxYB4ysHwayNXcMGXvAJ9R8R2fUapcVQP0qRVfZPY4/o1mKs/R6hA
rAQYImCUC9SUurIcAPlePSADpvztNy8VmMTwUaHsz4LA4JNc2BIZoOESkpqgpk3l4brSnyEjUnvr
LtWMahmAsTMaHRDxVK8wjDiTVM30K7M0w07b/lqHM1WkkzY5x0sB8+jXhchbqWcEI1gZwN4gjAfg
ZV9BU8EQ5tAsCsgxCctFrWooMfRC/WWldDRkJvXs1Npv3OqHKrh9VE9ueSkpdDBuY4Rt29I+mDWx
pcMwHOkX3PNqIhVTtLGf8s1Kp+VY0gZn8tX8QgWyhCqQG35XhxoHy1vtVjXDaHsVLP1t87dvxpR8
i+VZQfK6wowRhEg6gpM/fs9WCNLKnjSU4QofkqUqAxBCa6H/Rnd5fgIkoWFBqyajS8LKyBcKn2H+
+ewD7rOj0sHtjRhsZTO71fuqaeVORIxDP3bjU40Hx8yIawlw3oK5N5taN4qtfGU6Bgsuk7Sg1qxr
wCALIREMhmP3b6iq1bGmQRXrI/0bIH+S2eAEToGkNgbVSZWdak4NDN9z9uhPZTr8DTmTl8pDZhk+
xi4evXhRlXSZa/4fW7UVsHGXZZCPn0yYA5Vv+mkJQn4iwFs+KA+8mxdMubAUu3rkX6vmfchvVzyp
hOqrpVlKfVytQzgTqc2OJcPVMXyEvA0dL037vrgPZ8xwQ85YsY76CbhzR+nE05D4Yq/JuJ3CVedX
i+gml3HfvdXX6tghRxyRpCv6+0gJxjiGodKf0Xr1qYIe0wLFghQtlBVst8FvznIKgtZ70Bfk0riO
V8KqgQw6U6/RfAO8i283S6fnCQrtJGC3jT6Tpp/zAChXvygWmL9U4vhQ92Gm5j708Bi4FBXl8FWQ
k71KzV09GKy0yn3Y9DEA61sAL830mUGa/mZQSZm3siD7xZRf/HeQ4VqjXdXH1fgl/3tskxfVLICp
1HRK6jb21nYVf86UU4ec0TajdaFwWtwIMH+i+ohswDo8sjadCzgp05g8vz7/ogrrWcP2bsyC4+co
AQaY3eMPOHB7ce1CmHH2LB3TzXORbF6L9K1dLD9jPSyHIKLFR78jyELp+gTn9bl0X1dTpdbiyABz
Hgol6hRYBI64Fs/eebtj19GrcJ1GILpbTtqtbp8Nbs6Sdfm73LbDNZ80BXeJDBccak+yhVOOQgVn
5UvbeH+5f8LXycpN1qGcDYAdxVNUzQTjXbGWawukI0vfPb8/Y51G+bUWgKxtrAoRW6o1uV9deGmW
8o1SMhIci6JvyrqQmMLcGmECelmwXkcY18S5T7SDwStG3ZyPuKsjFBeCrOLmO7aO/0XOPsZeE63o
fWqhs77o6UJmJiJDUA8y9VL7WhPn2nyjBEJ+7/SRztgSpxLkrtsKxYtMW9S1cYCpZuo1nR9NSNfB
aViQZ6j7BQ13/I2Lbw7b39XlPc2eeZ3VJjjFt6dDrQy02mN8vbvn1kqap+iUCwA0s/69R5UppMDj
P21tiaEJbg+vF2E3++wNid73NMWPQ/JtDQ5XdpNtvJvAUzehO9qvm471wD2b1Axf4p34oN1Ddnug
mCpGzeVho7LUe58RZdjKoRgXEAQtZg23v5CXjt0U431uShB/mJtmNbDm4dMBF7hVj4L+X+L6dZpj
mvhdfzRJRf48nDTCpFwW9gHzgH2tKBGh6/8gtcMhmBq18+IudTmK6MD6a2gu0NzMi8hPZEA8ERcx
ejaGKxRQFYOlx9Lbd9C1iTt02d/GA+YcfYbCDmPDfYCXfFjlYGyMg7BzE/isly5sBr21gvd1eKK+
aJXmRtInC7HU/TpqotIU8OrYOXTv6/ViwT0H9rpPuQNckiFLsQ4UVCOI0BS8vjWzcqFwBnuZcBRb
tHF9UNwth26DaZVDxl89YSlNyEPKp9nTds1EdA/AWVIlaIC3kLcQoIjQ6cV4eJY0JRIm2PChaacr
FGC126imqboDE3NqKKgbyv6KBhJgBCL0VpV4oFCx4SLJYSjD9cQ/pzyu6hVjw1LN3199uCaqR111
tAionh91LC0wbKfuZiqFl70eaNR6lM1wwAOlf5TksuZADAocL311OzHjJ4kya9ZKGu/CNbra99Bz
HhEpYd0BBIFJYBxJMwcIl4L6kzRF2ZL4OHTf2EJ9ou/ibF2qs8MlUzy5AnVO7oTqTDqkL/Py/CYu
O7zdLKFJcW93WK3+XiVoD5tCYvGr8/szKKp7hTbLt43aTE+WROTErzp6UNGdVw4OEumTVOKQz+gK
iabL/RVaV3SNJz6ekWdjZmWoCKpAyvegYqdngoiBiKgk9czDy7aSmYIdPBbNVIgEq7o+t1XSp9jV
COUcmypqoskUsob2VcebDnIvsm4Ai5HseN9lbP2SOI9G0w/UKggn9ElI5vkZvf1X2tMP+okiociY
630q8FAn+X70u92IkW3KR1zn7NJkG4r3Cg+27hljI87wx+YkcgDHLSscEHwVm1r1DaQiuMTn8xaA
Vl/6kX+Tk60X+jprA+m7hVJNYxhu7xh2rV6afpWwI3hfGp6tTR4mF3ZicGUPzHVfNZaDCLPn1Mte
NAROdoUTHHjJVyNJEmGIJkl27bJoPovvOfGzi+77rRZSZoc65VKsxnO9n6kxfQsLJAkcjMWqE05s
Eq4ol2HLrySoV+IV8/BdHs+dB+5HZC87ZVjuOIsnqFfVFMU49bB4gscdLGtMQRFqQHXAM4MWc+u7
q/+ebJL+hPnVzVuLSwzhmXKi0obz4sqyunYvPkyclw3CeES7J0njI9fb1g7obzw3gwH6U1yMYrXx
treoW1NPPOnlCEUoK6/MARAsEV0WD2PHp8Vb6vf9vD5hfTknt0AZT0JcTD68C7mKMVm374jshDEh
snL0ZdoXkuTvkP5zcBQwPwrwoQ68e/0Fs8G0qy3yyjoVUvIz+EDpsHbXXHTUZVmj9py+ccvY1r9E
kQDjtoKXyb3bQEc4T8xEVqrHPsV+tKb4PXlYobOSLc0iGQEIrZJOcE1HasfRWWTWmymDZtP/7fyg
0fMIOUPIEzfkzTp1GkEIf4G7i7zsu+THKo4VRb/Ucu8iL0KlD7AFy3LKdcavw2FF2EhyRf4NGl4U
UztxymLZlAzxSQdjgElVyxYwJVvMOGAn9IU4cz6w/L3y2xMc+YEmdxoIBU3g62VDqotjWhM8S+eB
cE2alAtMe6lydgDIY6Pc6gPR2+cuZBNp/9FdGl64prjU0GIb8ZdaT5YgWE/hvCpmlwPuvcm307Xm
4RVyzBPGxYkMpRD/cfbtwIvOH2hwq+AlVmdPXuYdvPsyLaKlqU1baU/5pVhnadZBT0NN3vsJPdq+
HpxdUL3V+ySaaeJ+SjZkc22D1wWYAXMhl78fedB1amdjk1o9AGA9hIgFwzfXIHNBTbKlnCtCdLoI
ngZShCWrCLFRG2yscbKHCnTJBln7X2um4lWvuy9pQEnUo1Bu00wBeCLq2nZ/uPYIGcf1QJ7pVzj8
oN+LunJqxN2xQYlkZGcaVj0NxPukeqkHqUQ0PjJF1sRxNL9uUeOkuGdGRxlq7HW1z+Z1M/LuN9Ny
5649dBdR5J0cwJaaOBw+CxGCSMW3ZmHS4DrMmmoDokda07FxxwucMubBBaQr5eHYZnTrjvg8c6Pa
IWJwU4vhWvlQHRsO2FkT6ZJYtu36mEwbNEwGYzv9Yaz2xHwfa+d9V+uGwrb4HB3ygH185TsXy/DV
55wDdzTkcBXxU7OVgnnYq5l8w/85mWvWxs6Q4Z54oulLs9vrfeBLiDdLly0CK3NE765EvveOuQsV
cJXpArS90CNoslB4fQ6j/fTVBpEOzTP4TM3taZ5C41lScWCvA1PuttzMRFAugEecPWYaleCnxlCc
u7cG60/XtiQWNCNNnr8MwcLT1rkHJtl7aJxfnSHSnG8UexnV+Mx6XHyGVbFlZ4gNWtgGtr9BWOlV
lL+IEW6loF8B9J1jttPke/CluEmpM2NUZyxq2w5WiBXnL/JEhKoGl0820ROpcnzsr0+HKc75iGZw
/3GP4a+lS/ShOHv0N3bHWggLuAsdL4PwtXfk/EWcEnwfppCHS374orzQh+jNoCDnABLpEqI2nOQQ
mS9wM7IpCeQCoIeExO/XjTMcJrv3J+wMH30nmUMNLSXPBjIOtgq9qcvSs4PAuuYly0PWLlBfrPfa
wrQWSdLAJo/ggvd6YBYdvEQFSPmGFNufkdY2TPdpaX0jnbGGoh+izb9st7NThCPYx4sfF45PUQKW
LZft9O30a99RxU6yzlBHy7SFzmld57ZvUksTzLq1kQjdSMuSUBGwv5233t9SlcMHNw3uoDP4R3Fx
SjQPUTxz/a3r8nGx1o47N+H5WBOjVzZv8TyBjyHodQ8PotDh/PJY8vnsqXBxkkLMsQSG8zz3ZE5G
s80qgz2yFH5pWGMUKBf//mI6CJN/RbSTEDMrzMlu4iXPeKlHxAuUzM5NKCrIouSrAc9Ju2NwYP7R
qixIHAhIGc8wUHBw+22+ki9hP3Kb2e+flpbFxV7E9CxdvGae4IPrfmWyZ9FHr745jQn2POrle+Ec
kjRZiouZlIE2av1qv6/s66HL4CrGFj5BoA6NgaAvbwLAi0vxaT/E1v/U1pcr1DyF30HhtQ227FkB
gkG9MpfyCQFFqt2Evp863YTlPVxHGu6MitBfLi/deeMVg/QCWPi9n5D6IqkrGDkTs/uF/8KAMBaP
AjsdqESe2Qo7GzU2cfWMacrMrGm5R27tVl1KBqFJVwBRD3V1bpf85yUj5mPlhrrhvqKcw9Yjff6Q
94gwrKWORhoysF7pyoOeB1nX31d7PqWwPlB9g5PZJdbdaWO8JL/1C7Ag6u1cd7EkD114b4xa9gjB
/qAwqAqhJvXe3Qa+wvTexvrSQEE2t0nEM1qSIOyGcWaUU0O9IAc0rPpQ1+sqTXcLv14y1MXjtRQG
MznGuxcQeaFqtjJKwy2AYqdicYdbibnnxEL/aOFsqKbeBFGt2VVwNSlkpXgpYY40HhePpb0TiSyl
O5YK1jFZ/lBxPxgODqWdU/FSmvfAzBIXuts6TuISsfobaJTbiP3XcNXabUFt+TCy7xxO8qO4ifk5
31vtuW/P+EdaME67ByCvsvKCrpKxT/GWUcjS/Dejr00KdjLI8AxOl3aPhRZR+8fDpg3LcLr/ZOAW
30nrVwJwYr2RTql5YmTMx775pGw4pvmvaO3o2X1cDXxuZVWnIyfTCn3H42tMv2Hy2nY4CEjN0kD8
zosJFAghhvWpGCeqhSMT9QsChw9sfGyJbFqprdWSbLZsNHdqTZLaDMmB4vgYfiQMDq42UyH6mgoW
IBoXWIjEkLJISo9/tZKgnKDyCBEvFT9Al7SjgyAgV3VTcUh0kmEdUaupM7VFBIZVnvZPemgGPzic
TVyTFHmb/1hob3XksznJjE5Bn2wl0n3q3qaNj459xDEMIvGlUyIC8fGIgLpLh67K2MMJEOj8tO94
pVr70xAoHqlFGVLyM+YBzApVMOtlup2dsu9Wq50ng0040xeMY1431iUKphTppdXUIS/iP4fF2XPx
9Oo2VWX75Y1o5Th4ZOChc3wMBo4Q2M18BBRMhoQD6sa5gNtzYSLO2VJFknzqgm630qTwALfzeRIV
0Lm8TcndzYFZ653ROShw0TE7sSDMu9L1hnuYmr4L5hPbu5EX8JJJVhETYcN1bET9fFQdAn2Rjl+2
E0Ppa0L2Jek3DWnzq0pBIw00q+bBgV/QJQ5dhM8JPvbi8pqboFgKK4YlS1fmoTVTeU8y8jjhSMFF
V6mCoBF4Tpne5vIMozw7hEBsassNHBKX7NQ9UPuQldsXTbJQffF5r8m1LjkNo5KMFDj0V9oWLmFZ
SYmmB6ucp0yL/D42nBt7EiPXRy66nm6ONPvN148uG10iHz/+55gkMuAN397bxmUABdc2ceShOfuK
r9gq3IQ1KSt/sX/Bz2Kz4OdWXFkIYGsy1j7ftUZgcsNhEsd12ZHwW9cEhZ5wyan/h1aZOJ+7SDNb
Y3W/q5jKxkmvTAvGpUdaQxX7P1TDQ65YxoVWVrYodP0Kwu8T6mDGw5Tz2VPmvhWLME+GcKvsR+IM
Xw2QavChQj3F/2NWpT9i+IiOqOs6cgOpJShFfDbTnHHiUOSFjLAxq9/UEnqlh8mFT2I1m+mWBJjC
Op29p+u4wiZ2EHagEuMz22JGxna+aCin7XIkpWDF4hpqGrfJSDpclmHHyjJcU3ehTE72ZUtjtOL7
1wR8J3WIl8pi9gBhsz27agXiPYeC4cDh4agnk5BX7uzxWiH0/zM6UD7pjf9yrg1j0hRzt8Lc8O+9
ZL+j3LFUBrdXin6lkyAZeHeG14mcRrvgzaCvncq/Xk0A8JHG/0OqgaDPcAnhiG1KoMldwFEUmFSD
SdLLaJVbPLTfBuhapis8to7dHtjke0GFZIKKpi/Wf5+7Irqiqj1bVOGrMQ1eCE6UmU+s49GG4VUD
tW2KTruaJaCkfbh/w3sZxB3WGLpTVUFyx5zYXoNSvriZZ1NUPAWB3tPwyEt4MZb9SrolQcBj6pP8
tdTSES4FMm0jaFdKoU6fO/s2i2aqjPGM9EN6CinwKT8F6tKyHYaVMdtA4E4I5dStHUGI6/Jt5w4/
5xqsNbgt1eWkPg8+lVqw/Ft4c6ajNy6V+xz2D6IOwjpXVWquGxSZyBKOXffi5wk+euJdo8exlXsn
5vic5yav/KqRwEu1lPDzzRyCqKpc1J6JR87HYC6mUvaTN0NGM3NYt5/McS5/EuAQWpP9amuOURkU
V66x7sVGQT4d7mGDQIZjhaly/dAzjrJJVyfOUKCYodx29FwBIlHqjqNbt8ZyPzO7GeCzYHCiXQpC
+nhCYGnwzTi90d30ZasdIo9B/Kdx7NUwoi2suwjEuU5kwHi6EAnNYtMmCu5Ng53gNLVYlvEJQVqa
ApPLDAPQ2r3AqkK6FtD/ke0KYPfs5NUl1ZeHK+prxlNtaLBM9allZnkZ2zinaKvSCHsloJUoXHWy
3A0pZzocNUpJDLJNcOv7H2wNk9s6m7tpWSJ2CvjEcW78ofRmDpXnttikdV1j0qM3+VL34J8l2epQ
b/96CTIWC/15deaaSsdx+lPC9WUgRVGfetDhVTgbvKnR5i4SI2bTqNPavf2yXGwT39mixuPpZNt/
uRvtRHumjIPcL+JKVkGNntCHWw1oGBnK54WYFpwWDIrRmxX2EAIRA1iPw8ei0hLaAxBUvNqh0ECG
2D5ciX4OJCqHdRPShTVA0oqGsaMUaKoN6yYON4UkVx3s1Yo5mlQrRMSGevq1Z8rfbrM0vHeMAmEA
BH+49svsIdLb1b6UnkQo0rla9W6AVsUArlQbq5o5TUsVZL2GNoB8ZWoCWXri5TwvUuiS+3iSpEoB
0TPc3ymCH9aLIyxFSmlht2lg3DCVgnkT+mESOvZQL5WMUGKvO8Vx8sPnEYsIxfo+mgWy2Gn8kgSv
gH7JrMIQ+6CbwxHCZkLiRFJ0MkTl28I/I0ixnm9IfL3QG86F9AYQ37jqwhM57G0QW+zWMacWTlNj
tUgr6tR9RYHSydEp4cpmVpVPLQavBi7s2EKFI+HK4vLr1bZJyy0houPTcExJq8E0H73xwQl98j7R
Od9+LxN2Nvw9q7b740cD/HlxyAUUMBDB93DExa/leOuatpwaX5a2vluzUmH6H9nAYW+mQ5Bkm6Ip
8sHfdzmGx0D7hryfKeQI3SC+4DUUXCOSa3ob2DLyt8TEE4QdT/sUZwM4qhIIAqgFC7EVdH5E3Au3
Xkd+Ri9iE4yHgpQ7T0zEhkVz5iS4fh6L3Re4qwLgGG2kbPv1TXGS30xYqiLxjAjTj9hl7KBqxXbS
6NjPib+ubrVrYNQWdIgyIloJX84vn9L0XEQPHPD17x1Is2rxE6eraEyaJ8eE1JPLxVZ1dEct4lay
evimJgHIUr59x9fwq8tfWRtsEPVqt+oT2XEMJcc6HJQ1mt3x+LXzEnnoGPf7xlUQlP2+UrorQ0hg
y5Nng7eQ2XtoMaN42AhFJYegjTdFr7oaZiZG3sjaf165CkZkYD/N/GjdkZflDns2S2S8u3N6z2e0
Mclw85pX5Td/QPA1vTA6wROa4qQjcFL89dXDzyy7mBXRrOYqSz7pNUCR8cEeRMOzp+NlbkNnc3TB
45mvJQoT3YCH5o2or5h9TOXrgCeP/+RD+ueop6pFCDfWod0EDqa9k+nsweDtWREjoaDrEtUZL4mk
u6M00h07cViom/Z+JC6nEniHda2ZpsPp74bMP5BT4x1jzHsNKE5g4vVmH8XWp+zVNqpPMdOM2K3W
Nmli/jGh8ePrzvaYGsPRemhorm2rGX3Ry0Gm4YksAP6y8v3CHegg+eOsiHqeJ43Kt4zpfp0FL66u
zAeKkKiUlgfD6Wd0T5+XEe0ljGPJfFdT2Rs1pQ2lP4/i2Oyqlh9tVnW+hqSw97jrsymzx+msZ4YZ
1rzUuKM4Cbgbz7EnmDtgPCBOTn8MBW1/bqx7SUUCJKr64NNY0O8dWt0duZ+nlkYDyvsyiGuF6AUt
ykxjZeC/yFEbLgNYi7tLXvfk2Ng33g4SrbQFDNhnv7UcxiM6GtG3sFU1/cz06MpNQfj0gbHScxpA
hvOAXbRodkxO6VOcS+BGZ/7z5w57/IO1QwFhQwb1OIgf6i/Vp+oBwzymU6ApnNWC2bYnTHQIHnkb
P09Z2XgBPAg9MtIHNOSVLKECSpsyTIR/w/WRSFOPnlD6TuJ/NPRNScMxwENtYMguDvbwIOky+y1v
mCJOuW0+EXxwNpIvChwmP1TxStzbmRBqKRnYY3j4McnzSw/9bkvlw+EcVgyDdEJoYIAixnAWc3Po
K1cRacPSrL72uuNq/SlDULfsewBwzsFM15mn/GopiGTHD+cJou55o+pniv1bGFG5IjwFxKZKdSGg
SQwcSHV/16/MITPJ1mQdmRk0J0+ERozIoTyH0EOCiXq0i8WMuEyyqwAQqCMa/YViAmwRsGMS56F8
oYjwPQJEeOvkJSb6OK80zKaqxImNSRvO7xSsu95qLBaFz0oK+TK1c1TOJBNpXi4dtk80EYdYK449
13sRZHqZTHi4mZcl6JtdIQ3dbeYejU1Y4gvQtxhIOhSme2VeE3L2qX041E+SwE7BoKB5oOLPjfVx
FqzpdBHRUyS6fwwTs9q9piF+kPKYxol8/gnGugCbRmhrWtSlbLww81nOWI6r9bvX7d7jLXJSByDa
4DyAibKDq/oA/6m5oiWj0fbTkbvBYdjcMpiRT9StaPemTbZzSXgpapmok3kNJVZXltpOZwtCCvX+
97go0OPNuq5MOnu1Fw5hTVZmk2B5P13/tR0TbjxlkY5waqiC5TofK4aHFqE79Err+CQstOcPPgw6
HaakOkWQAvNMGIKujVeymZLlDmdMoMV3WR3/vdX7xpLik0O02r7cV7KDo5OpycYcdFKBflBNMmh3
IJa45BiLxJPw0zPdiWpceA4H5nWfcoa2a5R4wsZs2OjkkKoaSIu5nQyPZg9Fe41CtlG99fS2PMC5
kpHu/VEuDr5xNcb0ltV3pt7Zboc6ScM8nf3KeCWstFUoS8cdTHFFyNQKAroIoqON/L4NXRBJs2P5
VP/WDT6KhecfAyLeE5P0pJnpHH7ukVoTLyVTdGo0bA14rcTP7URcXIhG/vslp37nwTpnSGhAjaOa
ixH1aT6UtsHUyyGXUR2xn149YiIS1pWpdcu02jQt8LMsGYuATDDDJ1gwmmO7Bot1KgyKF3fc73u4
fmN5uB7Jf1gEuB5enBST9wqRwStX+PIBJTCbqsOLxfUYXkC75jBwHE0ue+By0RNQ1J8cl5ieDemb
hRtbuwPKYMW+CexozZGSmnPj4To3znF1ibt7ERO28Oc/LNgwN1TS7FOP6kgrrGo6lSYztySWc0UJ
P96Dj4xAslXjg1otNieaYByhZpa8KLgsygAKLldSXoIsrle3j4lXaLrLIYOJhhMgCQZ5Z2RAUzL5
+aQ6w4lFCxJeDTRwYCzATQV7tbEWfYRiVxJVI21A2rRrx+T+2el0hvDMIXyVy3L8AmSu5/Tp7ZtH
cWWR3bhEDIx0IkQbVhwQPoUFu3pyj9OljXzaQYhU3ArArnHeuRMbM2YCoPgtDdFOD+kAhksSNkoP
ASfSIUy5FbkFIhmcIlb+i/TLeow18mzpK2H9WHF9ixgbqPH7LmvOxrsL2mahQhhxojFGwhg7I0eV
REH76Iel5cX6W7aWzxSlld5DKpejoCF+/leU7QNo/Cg2vSLdGV6Jvzzj6gxwX5MHHSeUODtgUYro
ZRh4cEpzjaTJQEkyPoZSJ0xqk6Tk+Q6sxsnVxGPjOFnGthCAYdaXSRnyj2zcbnIRznO9CL6AsMQu
3ta7j10SGmBiQftp3OvFNTpBDXAePp0KDvaC+Whn2g1kRDij1F1veMfvl9GyjDKvvntpbkuLaR5D
U+/vGojx3QjK9vHtAA7fEM23UBbz11gucEAVGS70AKDaj1Hd8P3TGilYnqDBfVakJ7qGPxgg8CL0
NgJYO+gfKtRGvg7D7wkzYqGDDpcvf/GRhoS0tMU+nRibs9oN5l71aN//FvmuiwnVSwQQIkm5tfce
vmIEvGD1J3tourNZhLpH/+5CpDtkLtq7EzqXHjEEZxl+hJjj6onXFKYLGGnAgKnLOgD+EqsHoMna
XI5Sax0WVldOubmD3FZKiQc6RZe3VVtkBrqhHjtfQ7p45f9tMWYuwcQpzngKWdnS0UBasnD3Csx4
KJbHEanq8GzaB1pv7VIHW+bBdPeeREQVAQd+mPBcqncim57R/7woWJOsSsAKJcmFZ9zobVW1/lCJ
j37+MxinzXHaPYxsRlkooryXmFZvv8JN7f/YKn3vNfVZy5z1sXtkFJyG+1SMJsgria2vkIazE5Iq
5fSl0guncvJqFg7c158afLSupq9/LB14y2r029ZKJvltfPQ4r12FaZksxHGE8eEKg8AKNwcRZA28
2dxQe0LekhQpezv9YuEa6mV0LQuDBBFaa3/5QMux0HgjTR3zlYyz7mFZdfQHcuru7vJZUHGLZzDf
Ytz/F1RBeJHHB/lX4ePur2wMI7CVU4PUDXmYA4NZdG02MLr0Ha/dBzjx//uoPnZnOklKTWpeS9VH
9EfaPX/oYZY3g0KRzDbF1hdUe2xgFYoPdSU14Xi9SAMGswsmBreovn8EadgAnntXu4BswCvX1MeY
LQnL7wtcFDPvptW1WENnufc+tj0GAyLIscJJv/LtIYZOq0bMkE0V0XGMHQAMAoPDZz1U7jXQuaB2
XEg8ko53Qp79TGCMHB8ZCTz5uiqouLMrIew3wjWv0eEfl8I4piq81dlYS5OJSD7jBFDiUelDAsq2
1HszucHEm12SW0YBgx3c0jBAKxSafEoZYbtA+CijPaTOx38UyRXEVGWBiF2Koz6st9BR0oeO8Xki
mBW0PdGSGjf0emiSCK03RbbIdLKd3GY4ZEsQNbCc3OZzrSFKCuAzrhik1QAcxVYUGyNT3Vx3u6dc
fAWT0wetME5MOtqTgVuwgsphrtBTH+0Ydq7TDGfF46t2jaEPlsvdrnDLgrqXBw5yWKzcOJO5vl+f
WrQjgSindslIQ33wIXhlTIwVURzEC/6ihnE3F7ytEKiEJgW8MHymt3US1AtgetyOAFz7rlUZGd8A
hXPJfiLFzgnJRR7M6A1m3b9xlJNupCceRWNDqsrK341+6QWwVg22lrYhtunN6zotaFkBdHdMSUzB
WzgPfZmiSayF/ClDj3adPHE+cdQHl5lyUC4NvspzO0FeLW0Au3bf1jRvNKP2QzaPYZ0zFQ25fWGU
zUpopb08CtJddmZ4lmi+fSQ902ZW3OYQOOVb/rslRZVuPqU63yKUSGSMklScU8aQcr5QXLdHwe9q
Uv6CSoBMVE77DmU426Gb+cX+GWLaUR4527xSlZmn7XADda7VWC9GZUsph+K7eaofFV9SzcZ8gSvJ
hS8elaLZ4Hgk6EShvcnGcnUQRw06L+qEHgVHudut6RCO8JygquHXkAS63FeP8NQvwU6Ll8FqjsIJ
9nd8+j1FBVGO4mOhWl7Y+Mc5lYFLxHHbtSxBBIjA9jjyovL2YFkTqDg2AG6LcTdaC5+5eZN+dOPL
yzLpjQlcnMLB+CsX9HvGP4QMprvgXSkpS4kIpYZVuOzvYDAh+N2PeOV4hJgR9TSlDCPvpni3T/o5
1OZQr4Q8s5yY2BL5XEejhJCc4V1u1WfWUfp1S/wmfUBjZ0AIJW/S5jVMow3baGisqnXXhi52570w
qqKGkWdPamkQdOVUTevITNcCZJPVL1bcbQyWkVdnAd8vVUQG38tVB8MNmqsqB8LC1BszeU2uyqU7
IyD74OZFR9eZ/V7BH1xI290/RNzHanGJ906I7uEqAkd+aJPKmWJ/Oq18R3HVtfm5dhuQ3MLSl8qs
DafgnGd6okmpXvpSfyZfuigc3UaZIXLJQsgCMHJSYf1R98RZyZBeQ1Aum7YVW4WyuxvZKwOh2u/g
6OEvx5K7C0tbsO9hoOboiVjR1H6f5akmcnlLecfo3g8YP6hQg+Yk+N/+ph5UuVvJy3vyHUkeCJ/+
D9MVnAF5dl9TkwN6gHib3OI1YrM/6qPmsWoNkRqvMDqDZ9I3nMjn3pNzGj9cO8GTUfl2GpZoLqij
ZCWXNidmcwNFXsM+02+uwa0NbrMC4LuNDfe227b/C0JW9+LsQ2EzmiYNdCBj6iZvUSwK1FHZadGy
PPGgfAehcWibi9D5AYqVS1cKemlogP6LvnYEGmhuGOTCc67+ZNWyG9tPPW0lQT8WbYxLasSaodYE
qQqmRbNZ/A3IYBBpWpWElOncPbwgFVu9L3O9yObN4zxhszEZqxQAJG+lCPtGbFu6vMrBMLu+TT+k
gU7ZouH6nPu1tlOpz9lY9p4hyjjBzR+GTPtNei8vhj8JcHJTOrviCXVkUHYFkkLPRGt+GCbKaNlg
2Rv+N8GdiOlmlAlt4uZxmk9wMFWFDeEiVBM9mj5BgBvqgc8eKTMCjnaJOOVHL4ptNR7I2nzoDJJX
sZ37pBB6VV9WjGO8lsyXJOlZCHicgK/7ICf034npIWukl8lEWz0TgawKC2CRvnWdYLX8aW97vEi/
r8dNzqGGkBQxMiZUKLXddePF87s0Mp3I/z5kkSOWAebNK2EpG/KaArYsOpy0CDNdFZnGQ9cKYt3l
sAN5tkBx2or/xSWenNQl3FR6NcXwWZvSGayfcJ72Nhg1YddMEel/JYUCAMVRQMZpvgSNfvh3/bq/
0tFOzyN+bjLv0bNXoOh4Z9bgS+zfYEHV3YoruMtKFvZM9fnszgbLTxi/rwL8zHeyW1+dc5qP3feG
xMN9UzJ9ESrjanmdepJieppvJEc4aLJRLMNsN86s5qEPxvu04KjE74JqGaval0FRrsC/dbQ+Giz3
Ba3acW5sA1Nr6ewo+uc8p1qUIX/0OiWkTyyzVpXkx5O0KfcLP8C1uaU7k6zz66VlRqQ3I9vUvhkC
XM8kTHq/YaeaXcXn0e6rS/T35nlzEnC1eyvClJgHouyFJ3HwAVuoDd8DO5GOfScltVFUghA7L4au
e33tSUq6XGzhYX+pIg1x9ZOE4U9P8ipUgg1ODjusJMCa7OV/j24R2Cpr2XragLgsi7v5nnKQWEL3
5HvKq+NhjbZOTs4lwJVDhzACnnttgrWmqvuuhef+6R61/spp0R63LqiHltXj9OCnVlx/gRBXGtNB
gFqwUvjSUO8wCzgbBpIoh6n+4tfgGcEx5AAriq6ngikd04IwgkqjeGf2XrBH0VnFsWFPE2POhBYF
5t6rm1uWfF1QfPdPDYY8PL1Z8Al6FRDbmjGQA8gTF5PHK6bWp9OPRylBlviPLSXU7MdvseAAaI6j
iqvBDfklw4snFXV4ATHBbWcXPkjYPXLTArdyY17q/hyAFDG/RuYdznDrhASI8TPrfbN0XR2s4JV1
SlHc2pQn6es0j+6U9lpsCTFfOAEpsPemuDJBOvnvWi+RU669mQ5Iiy3JvQtM9RrUxNvxjzggmW7o
eYfvhYSqwGTJOC5x3ig77grUOO+6pbRJ1sTtYL67kVq/FJ3ByKchEMZrGZYldmlp7YruDWiqqCPr
gCpLLvWs/B7Hs7xlAqLyT29TfOXD2cISQHt/zv2gMMqyh4yJAGV9TS9WmdG5qf3OTwxwtjkBJJx5
IlNU4I4R0wQU/KtrY986/SV7iLhv2vJqFD/cZgCDD+U+9CxPHVuZC0OnzD5dz8gqREm4ksX/y4na
JTpPyljW5/KrhFmVIGdEfdzRsNx5v0YsWUxAquRs15HUx0BJcKG/G/RAHX/Lynb5UkuAoFtp2Ny/
39OJct2UDfYK5MFmbk8GMGr+1xS5KTYcD/SX2TklzB6PcSm8aoI+smyDdihPEKANQNwAXjah37Ji
RWhPK0gyhxIq+2hSFnGIs5vsUj/hiUZLwS+zgfmFYX9WYgCKmiINZEcjyuf1vGtOWJxYtmLoqUlv
1IZ+1hX5wZu8pbhzE/ZoeQtFfZ/LIKqz2U9ztzQ/MwvaZ8My+w94cttrWSG7SF8fH7FL9ByOO1tD
XCm7UgEvqrLUM6qLQAVoLDWINU2gRAYgPciHuOZptazMg2QRr8l+sT8Oq3AN2hrflbBr/SwP4jdb
xQBFcoS+Mv37W9VMqDGqVnRnHzC/kAi9u0DR8cQzYb7qJdFHkKA01q2nC/X6YhUzdEolfH8wnpXa
L/s4H2sLDT94ipG4cZp8cmFv4ya0p9B1ISCeRbHpttlogYv3eGZeYpTOtoM3ixbbRtxXGtKIohnM
dglBxqp0sMvzztEuymb0xWRePEXbpd0u2h84f1MwInPIP8Fj7L4fYZzbX4CuMSzwpoRwTpyHdr+F
ogOL6ktWe+z/VmUWntXTjIyxJFA/5DDw5AsIinFKZGeD4q/jNLk781KnfcAGgMZpJYuKET6+3MH+
z4rOqwwmAsQqyaujpmd+l4hAi++x6HRuKoAPZoimN8uxKwC6dADk/VPePu8hdQp8wYhwhs3BqmAN
HA6/xa4c/ClxtNIKUhMkAGbxU8iUFM6NH9i/TEOq4qhsteuIsDd08hmS+w4naOssM3njfjvpy6ai
GCLw2gdLLVjV6AwTKJxqQJhIAGLIeI1rdxqQe4WDGB+kJXpLf4hYZC2SnnLjJz4G4JbV8y6e9kxs
H0htQfbilSLjlw9NxuW7mLZgy84oO2M5Vz7NKyTngZEVv910i9OgIPCWsEKaGnNd3RoDVCM7MfA9
BDb1ZNifFoGy9HFPWulPFHCXseeAIU9qq6CBklbPF5h6Kq9IjQ2WR7GbHyeez5yuT5Xc2IBxWg+w
3K5T8Lrnc7wbPME6iHMzgaujkjov7IPDIjsTzx09mnSERt2Mc47XhtqgcJL+tx6OiWAwYu7AR2QY
+AK3jt7DuiuGHhQyW0M6Y1p5lndwTXWtlHWA1E34E6BlbbxTcr4hhTs/feEf0WkIS2OQdwbt3zw+
pQ+clwQ9W6ZKxqrasOHpH2Nf58hpj7Y9F9RCDCJPuKK4rjKko1svIAB2UJ3ppq/dNQ3M/MB54TMN
qffxDL/IRjnSCJW6FdmYM+HmLI+OEKRsNZckBHT01uJZvrGpnxtUHVTyY04jTSH9nNCl7xs27VTb
JG9kZuPQtHgqsXCFENWPEmDumStfApaxik44g1Mt4QFzl8H0ibcBE6XDTMDmPScj8IQFZ3O+bW0s
I2tC92TRdINO8bXfYYClkyPUiTdGI44yCh/FPgxFDVBOiqeryf/KAWxA5dpwtIc2iGc1DL+Mfp43
qpUmOCyq4z+Y0jJEG9QlysSOGYNPZX/4vMliRltpH2nzs0PHLbbIrUSlhF8OQCLzSyB5Wk8IYLpt
pfxxfo3Ev6pUrVM3aGvkvsiINTK//oH1lqnEjCKY2K5kN4GG9Xp3rXFTpd9606LKSRvPjof5yzsV
zsDb411QTvhuGwYW9f168QQTr8I9yDkxE4j3Aguu+ZShqg6V9G7BfTlUcRDnDcfCS4FA0gUZct6u
W3LB5FegFhv35s5gluMI3NY/AoYcolklXIlAMyPrCTM8AxmxwYmszCo7avELCo8jM9wQvYWwwiKN
0B61EzS9ln2HBij6hfYC9BAJJGLlWQy+We1JhWYF2a+0E2eZbcNYGDQAG3yY6P65LChVg1xuqT35
72DxPnptt81lTZyaYBkiR1SiehPNeFhp+3TLoH507owYuhQW7NBt2NLaPIYKeM5Aj9WGOV3RG1sw
ZhpQvsqkAkkkbWVdLRBDxgcT+dIIru+//F7r0rQfaaKHxGiHxttO04bGfJRWEvNwnN+zMVD0mqrI
CTJB2QDdnrHZNVQKjddx3SzWkhCRZQjeB28x/zXIGt9SjQN/lu0RxWJU1pacTTKddQwfTiCl/9lg
LpHlZrs5qfn1itdqRMI3Molol1oTyLxbCoBs/KH3IIUwJjwM0opv6X0RMcPYqWqMprIWAEXLkFcK
Eh7LWjhRseL9o1gs4Mlsi9gnJ0W2ViaBMmEdqWm/WKtHPEOxn/nbGfnjPoHL05hx7InOYUFhMObf
vNBAbPY1URP8/16KvStEX4vnU9kCWWQGDWC9JIG3K/7xd6tbm8o3uxu0ryKwKDpeanAtzeitYL9o
HdOT2DQVTV68muy9/J2NxAZgXFCC3UayWI0pCYk69XesSjfBbJAoOAd8kLI891vKJo/IkOKD9bVr
qEGOiaPGbylfCik1brJhftLliaDQnnfgnvPhfb39zTMly/eS3BN2kuPETihu0hJRW20+3cG9BKh1
8/xO8CxyqNM+lWMs1OMV3khcQrxf26GKvrsh1NcuMpzG8AK2dDLEYnjXkFylmn5OwSvY/qI1e2Px
h+5h22fLQuivCyccOFwYVb1eByRWS8JYSWQ6mSMicX30X/03SPxog9oQxvdqPjlpb/6yYO8TaCcR
qBOrMfHJI4vm4VXHJqp9PDyizo87q0wRUz8rvdnyACpZlNbgpOUtoiGrxh43YxTjU9dXy3adj/DK
G1S9p9ui4wUrBYSwUmhrfTv1q8mXySVolqiC/JeeK4ELkOUkIF/Kz3adIFIwyCFEcmtjwRF54kEf
RCCYmpNQfg5SjfRvkj5JqsQuogWQEYl/gHNq2quQzlE5Lw11RHvjeOlcELt8E03KcSykE2S9Wh2Q
Abj8V3ccxgWlzrd4tgeYt+nwZ8hCVx9m0kT15bFPvmwlSmJhcZ/Gbh7/5P3j9xkhp7mJ+wbZkGh3
XDoo3Og0/GU6vlIzoIrArjXGynnyJzjg1doJhiVkWTPhslAimWxt0NbDfCghAUyBvy/bgaf81/ks
NIHXRQX/jCdoFwVFuPCWO2pMX9gNYewnSK59/+qVbni+pF/y/Oxe9B1oBghQcEVZbzijDozLYRz8
4EtT85ECgLo/2375T/ZS6ua+8Nup4DVALdibjj46s+co+It+XbkjcqApmxPf1YIQyFl/3zDHkD+O
36Qg12LUwV3XCyhB1X/K4Km/gufba0cIcYT9kEUizoffwbCc5lTOCJbAE3q527+cokejKK532exu
0f109fZuhzmscZ5v7zDW159iOPdspQqpOQJCqzSyiHQIGIeY2W9m+nW3CStC4A9LJR7lFbxziLMN
RF6pAnDGNx+EDQ7Id5GDnMvIhT4YQqLUTJdC+uObl0Byx+5ut+tBvOrBu44INE5Meky2PJ01Q6KW
y09R/rgptntxXN953SLaPRhiJNxtRu2O0wMY7s2mgWCYELMCDoUf+STkrC71k1gCWN7PaBKTUg4A
Q+oafA4nbltIytDlDuR19Drzyr7lgBoGG/aaNvJXANJLNpZnzRv/nVEcxaRbL8A4khLArUBp/wSL
Og2S25/Da3YPhuQkRyOAmNBHHGn8tmjLOfqVYvHkIBUlurhB60P7u7XrXvM6tmADI37j9YERPgvF
xLlN/VVoLY0FaqvnVaKxGy/+Yiu/QOt0o5vf3HMPzISrF1rLIozXe2ktqSyCl1819vmcJosMCYtP
it2+Yy+BKd5UHOp5C+PMeFG5Vw5KKm8TaxCnJy2JkugsKal9rIWa8kIB2920mVvDwE8+JUofEwcj
Sjzbn3uOB6xXyl98B1Fca8ZSPO3Ot0t3a9qcpRNKtlU9JVPh0tVOuOAyJ7QhHiUUt7P5ktv+WoOq
GR01OIoHsXFLslV/H2IzFfE8X5XHV98bJpP0siagoEUFOaPZS+sio/49MC586vTqcqFMmQbhig/1
X+drXV5vqdqfWyuq+CU2QyRXvVWwh37aLO/XVLNmxMk03Hgrr7fYh2AXoi35Vtu1vJzLa/Bfl6kF
iprOPcbGVAQNqevaoLUsvLA3HCJAGx+ZpNYx7aqdxkHKxOLUjpjIZcxhJw6H0iUV4LizxWDf42if
7AvWjc+z8zWc1nB8x+LXXu/IEg8U5s43HMjHxfnhwlsBbnFfIILiWhmvPzDI3czAylDOKkfL500/
3o2fgSiYPe5E+a7YzqwgndWYro/U4HF/DfCG1W4+YweuXBN5cMK/nRli6X3dM1b9p6yg9WcPq/cm
yRwgKuAcIa6dsZVJAX7tMmQwjqH6I1C++jic3uFahYWExZT8GMHOyOMsaggcp22E0+bFKnxa6D+W
5IEM2+fkpCL8PN1qGbAJyLaaaLr0A6Wt7pdRms1R4DpFfNl1s0HdMpJ5D8zgSL+bX4PZGRtTWgT2
M6JHB+auXNFJsto1K3mWYa8UuaQopS+cSiwU78AuEIj4xtmi6KPBwIFhJqp4BqEVlm1nHk/fRcJT
0P46uX0wkobJFEdXMVp14xRwUjCH9iZww6wgbYR6rXCPP8nyiqo2RLM5UNHaci4eUOhD6enV/VoX
fgqLvCJ/215UZdaFv9rMgh/XUD6EaTGdjPuuusk9/8KpfMkLdoeX1fE37Lz4iT9QqsbyBle0eowJ
M90ofmYR1gjYU9iH0fE3rhMTs1cFrKSQ+ljxW++c32Ep+mBQCVmFpzUNtBpZPDx8KkWiufKAm4SI
hPVZSvL+5PURTNrwMcvgCZwpHDSUnzJSlnyIS1OslGvedASPpRanXYOQNEr8aedkdBOtyaLF1PMj
ITd24aaOPzfXSVlN7k8yks66Kmrqen5/Mn9ulypByYxT2mkCEHjAB+2AIG1xSvq7OwQTLPXTZx57
dnzbnIT0bteMpFR022yClsJ6c4O9WM3ZHwBEm8qoUB+36ZDi7RCtdYqBqqOUok/voQk+Pg127YRl
X8y/ueTo4KOLv7UjX1u172sPBd19e7vqvFPqmZiy7FrPMewtBxHpglY62F4udQnnKDpzkqua41+/
sk1JMUIU30za4aPf7b+TI++zTjoVqQwaM0Z/VzwBO6++L0UEwbYpDYfp5jTYlFrnBc4Sdz2MIQwE
EwPzqGJueQ+NGXjPqr6M17fcnSe9gGi0yZPGnrRVF72Pmpp1TiQ2pXVkz0be5jOYc7qy2+qOAfpl
5ZrkAmgbpvjuernn4G48TCeLYXD4HlPjtJ6AhKWzMTXzrVLKg1ETHEP4ayuM7LPlqBTzCqC+K9CG
MY0qIRpKtqtgjo2TF2wE2vydk/+5jh3NR0ecnha36snONlRLuF9l+XFfsqOyaVsxoqbgNI8fXlrb
iLfzHajQERT+n0G0P9HQ0aR8BGAfycb0MYtU83jOSTNZ0+F2ECRWPpn3oFaUrHGhijHGyiL99bxG
F4NGeYTz5drTJXkcLgyIpXf8hr41QKP2tIktwcXC4bmuVwv92F1wC1FcDWbQpvJzgaRtYrKAYW1d
DMOxHmmo0NW+TQmhag3MANxoNbAn1whC/jfRPWjQHfvo50wW9pdO+VzVI20wR9vrm3lVRs7v2YkO
JVPHdykTtBJ82pbFteyRUkPTwUR65QTU2MwGqTxTmq+ze0JpUT7V7PHGMS30LFzKsMuPEkkr8rX0
QYmc06TSkcvI66HeNVz5/Z5tQsdur+E4JPInNmAA9cKcA+gFQfLs9XPRUOuCRJM295iK0F2Z+AII
2ki8mHpk5SXBFsJfYsxhaOxy1ZqD+i95ACvS5u/GPvDk3rAxl28cxro4ZKVtm8IOMw6PNunIQUtK
9sWm3Q18/6MSKP/zUIS81IlWu14ukzyvEPMZS/sXtaqjkfkBnQn40WrOpTHAOEB6NIibBXeGUTaf
NiQjaNrST+AgTEqm3arZBThJ55bcrNpSQCiy2uXEJvkm3prq6A7D8o0D0oqcCqQu+xNnq1COmB0h
9RAEUz7p6N3IqkOgWr3ItEHNGXZUFo7RrI6A18uAKKBF4aUTPr6U/MwZGEnRJoG1IkOr2hmiMBYA
9OMZvBP8qhnde6jxr/rVKNAwzW1HUXbJYWrViO10OY2MU/e1G5jY/TRpnLwZyDotmVnzWrhHq78Z
GK8yhk6aC1CxvTeU2lxqrs9SdiKmt4ZHS3sVZmH5/qRhXYZBO4LxS+ZJ41RaNwoswVIe8+uaR0/J
ZzFs8sZjH0dNnyLYPa4dUukRUA0HlquybAsFKR1+LD5TB2We9qap8aThlXWLbc1frneN+1amzg/b
wCLtN2EH24Zx0pIlOqWPoMxw872sUo8pq79/DMT7sRf2HWmRjve8ixo+lQ3u/H0PEs8ILy0/Un7R
DqYclMgBjCp50EirDCSPODmf7hykJwPNbnPh1i9c1A9ho+V2hTSlWOe2CJvsRXQVwCd32PX5Sok4
S/shJZVeoNkUyxcCfOeoXGb28eQdmIApM8El+SRDfnG/O4bBfyqlnGlLIBHheZX9ZJRp6ASJl7KC
9i+B02CCfuXm0wxinxFTFB0aPHXdHzdWMFerihtllZcEHWcRDwr8BNURMrq6CMhUr/SQsEU041EQ
Fs3wuWHYMJUrSWAknjOIS4IfF1SS+ZRdJ7S/1c0eehqT/DvrfZXO+k+GWmZ9Cmm57k70DunwHNKN
cm1/4UmMTV9t5OZBLWlJQFroRBR2OzqpBkldj6mwNhnFxuIX+ESBdxyzUTMzcc5DHW5nfgA+zPm3
LvlBOsMyFlD3T8lZcsJoL0cWZmfUJ3meqThPphzbVw2fMjDUlqFj/sMEbT6ttGcIVdYM1eqxWMHO
IoOIDNF7iXbgj/TAXqAwK7jO5BZf01cII/K/P3AF3Xw8oXt/KnPtc+AO0f7damMGZy7+Y4CmJ7jp
DSmi0q45SA9Tfy8wbHzu84STz6Cy4EXX1p/WNJ0eTvn2JsKLBcQ2JQ4+2/uIOCHKjJwO3j8CU+Nu
SaISyPlr/cJv9CuxNVGT/pt45be5xa84gBSSQYQQ0x2DvRhKPpc5iRCRUsn4CM26Xgo+tbt4U6nM
fXCeVFKupebzw8er1fQH7dgAYB3paBQXD9srMj2Hr7NVnLMFkafoASNt0cYmd25XzXxJ0jb9ycRY
Ct2Gz0JFyWDKSnVAzMNfy90Vq1BbkDfRGrYd5NR94KEzxw/aazhyZsLR5RfaCTEZNWm+2Tqfx/iF
ggXdIRO/+U5YQU7+bXDM/gVh5U0qSMXQUxS7s9LYEMTqDMh7e2N/uzJMOhxQG26OIfWhFqiBoeDM
mnlZH8u+39soypZHNMyE9Q/tQa6k/fBXHyyV9yF6bqzogxDBFue+2zN8HYUSsbOvRXICkhsm4TcA
brjyYemksITeAnh1SsWmYPTX2t6a4eEJzu41G3JjS2i9JvV6H2p7j/dUDYuCR+pSSicLZnpylB3X
nKC8zTNHxtCc74WiFDn9PvtH9S0d+yNgpkfg1J7L2LqSdMPK69Xt+s/HoibS1MqFxghc9KGBJlu7
zLH9KEhRpIOySqDe1yP8+pjHaj9phNXkhtfUZLCLnyNSaTzwyql40b+6QunQJyiO5btdcS2n6sVI
pT3HIXV0gID35ZPlELxxkvoBYlbzLTlkXOvipiKmJbQ0Y+l+opyaSu+Q1gg46k+hGsmZZzzjS7EJ
F6X/pFC88equ1HrlDk4JzqwErS3fbFHqL0Ec4A89a7ruZSynJ9X6jw2nxVtMicMO2a6Da4wDwMOa
vhWlt/IG+g2boHAXtuHXJ3uka//5rNhkLOFPrWtaelONCjhXxiHqhQsUlBzyn6IBoZnT4YJYpkLk
YKb5zCc3NCg5uCcA0Vx5IMQzBQhz/OPwr9VmcoRo34+3SgYO9kLanMrbBJ0QMGm377iFgq5UbJQ3
sykDe9l5oi4xejbTikrDoV4+gN87iA9tbGAIh2GizZrek7zwOX82SM0UifRRXsJlvN6HFGDLr3MH
Ku628QG2H8I3RvL1LbNZ1i4lvvWWIh3lBaXd6PMKxOeA7qfnJLiikZwrX+tmzgxD6mWEG9dNsvmw
C99WaDJLX9I72e4XIuqBqqThDTuqsN80lsljwnwb+T9qHsDPk3HqB8RvYi2R4zvF2yZ3K7ecsq5Z
Yg9+kz1ujkILStWjGYdCtSDqYH7nMKR9bsJKSjnP03djB+gnb0FHn/2I1msFqsucl1mN5VfEo5M4
+h6Hun5f+vRSlZT13uW06H6tVxHuQA0hKRwWC7vZY9nL8xqnBizQeMHRCP0tah6CnCiHrUlVtIML
3ReGM4iEwTwnL2QIIv90S5GzcWGEQuOkufmWltbZIGvm5u57D9PsJQvi4EAcYjT1+T1DQhKqIjFQ
lfqFDzUGdG9ZZZdXHS9yctdfpmt85FHYjyIHhue6o8W6IJH/f+38ndXPHt9V8gY/5Nsd4Tz1+mmM
7rdyZBL8DxvD5DsuqEyrdADbbz/TMwOLAs37qkDtKbEIUQNIdfrKb+LFdQuObV33dniBiYYe6Of4
N2pCf+GlRjl15Sa9syt8MDRcv0AJ937Zj4z3ja7XVRQYbVbl9wvRJ8d+/qbCsQolPKzcpsTKKZl2
9mWsXZp075uNzxdr4W6Hmw4rm7ZlI46dHdmzVlr/qiMCGalnRWkWgtC+6v/7npqRVnWRH6bv06C9
OcXXdxa6rpkMG2ZyRTwdaOQj5ESJBsTlF8UaEHa+RmAeGteEK/QSA65sss6Qym6Vxmgknwr2rHY4
OJPNgdvH2/YP3ULa9LsKSloU9Chx0uY1xUElH5i8LGbi41m7lL5Rxmt2qrhr7334UGyYk5LNUqhr
TyIGq5X+dQQXic/9ORu5Udblc10Z9jShpdVx7Xop/KB3vN9IqulfTdiNQToq1iVCp6hWUKB6IUQ2
OotgWx/MQeYV5YqQBzKdIYP4buiRHGf3RPdmjXVHa6Zlv01Kc4MeNrMc4YEG9gJuva5cgLsz/Zry
qrDvsSwsH/94XAcKiUHFH4H1aewrEkjsjUVnmkkH392XOqf9EnwYdvOk0/AGeM/CHIV19Z2uJn/p
fYOMOqGnu/0HUeGs0EuPwmgRyfSesnafNdA8efz6hIYGQ7P0vmizbEBkGtur9TQ/NU2BzqD0FENT
CbdNrqZulUMiAS5ha5DhNDNFn+BP1XDh/lG8wSGofXldKPTqvkx9+YI7ez8iHqIjC0gOnkXv/Rr3
tzvrfq1Kjy/nPySObcmWNyAe/W4GE7Mg9G2rCnkQaNvh56szG+C6taZ9cce9mihUbTIOeyEPek+x
zjPyOd3FxSIxNqg1GXBd1mm2zGaf+b4GUPBWjsP/nKmdhRs8ghuBtzEIwDrrbB4OoPJNI5S9fZue
jxL3wAZWrrKTnO4EyUfdEMsZtYzfNW0FtWJt3hQSOGyQ7Qra3dOUEQsIk3S5TbAK8L0+2UDNf2SG
r2Q6dyFZAN9yLcDTmNMtQgQQ3fXvR0hCI31lfbvkHJvBblUC24+2ciiJIzgg/rB4UO25vD96CoKR
EfIsbl5RAnN0x6tLiE9MS/eTrIc9xCq6Oyxno3qEAY6IFCQAyY8pNHWwAjmAkWTRf/ouCUyevFxz
jybDZHYGzJBTZoKnG/QF97qC5x0nAu8VGASSdvoBVWNcK93OvNfCd78diQK1BXt0jZttGq/XNiJd
JfXFbexlT+ltSlBUEYtsVIiCWDY19XcoNOlobRXFNnZGkpEciJW9aRzO2sWQ3FxB+sxqoBRQsP87
Nf6zNoG+s5vOxP/0ELiwY1sFf84qQ8frO8efTNhDOIy3L6OWK2vamBFf3QikJ10wCvma1Nphxbop
JU4HJ3OZkJuX/z3gloqA1osDh3Qi33oL9j4qgLyrM7EoIDRz+7SHTzKyJJtwLdTMPcdirby0mQUB
t4603lPJk7s20q1duX3e9BupXeANon6x/n5ltKxWeFVOxXBDkA7ZEMFYLuOVEWVFVpegx3OPoB53
3uvvx4F1ZwjPA/Igh70DgMJA7OlANSrKuLiyNXpYiRwqT+nRJgwmEMAuchFl8tq82h7ShXZueP/r
FWwxkO2eEHF7IZOifX8wHkOZcB4oOfhai6c9oxOAS9xbpG6ojKwmR52SFdzAMKvcrt4fZVPPKsdW
M7uy1Cx57KeDGks5k1lFXJ0D3OeKFp4/n1FrBp+cDxDwALFhxlfbv+Ur1+YG5jDwL+DA0C4MzcCA
yN2SUdXEGusZVMxqeGXcmrZ55EyA4rvE3UtH1DkeS7b59XrSEmx64sEz0Ku1Ijc1RJ28e2Jb43+d
ktKxRPGQCWHEgPlgO8/iNqkJsFgj2NWKX5SI66DXCpOdwbCDDpYfr2EL1AxLJY7/pR0CAnOC80hh
aZ2AQvFsBk1S5EBbu3HiwhTqFsNJhkCw7PERZtj6d2m+bb4YgkpInvnp6oOazxqw37jsBDIF5cBB
y+SW/ZUJMUyB7wTti4Jn1Bufcg7BohQbaUK2xIZ6co5U1SPC6kt0XYf36/EV38MnwIHdqGcPJ6w/
TzvTIpy/ZgZaz224iApXAF11WH5LNntbTsGQ7nnMCz+PpDgtcwqXAHHE/S4mMpwXOum6i1K584eC
a3RRrfhjtyX0pCgUgk+APXLBy+l073cISh2HU7r7D1Abu6I5WU2tUaMY2cVW6cDQDwRwCYc65VmV
s/xik0uQrCQQnlgjM2EC7tIQJ8xRsqEzVw+soNxJ2/3M3XEVHHd47qo+LDjsgYSYdeDL/pbbPnz7
3ztMqnakSuwc5V+Scl+gLf2CPBPNEyg74kq7mkYaYY7aEOEro0Et+RaluktizPfm1ifdM+twVgg0
K3s2mf4dXw7Pmx8M705kWfoC3pXn3x1sxPWLv7p4VEVUa8DFWW6TIm08M3bUQSAkYX2RKdTjc/PM
mA2io6dLSrn1Qr8w3y2mXpQ5SgbrdGvp8SqVdmMkZyw6AaIep+NM5/b2XloMLBRN8W8mq/IWANqO
tGLbaPprjSobJPEwpjMg+SbP6gxWxSRiAsU4nIakKbByHX9PkqB4HRkQLGjdggxtWdZM2UlxBMe+
eg9I+AfQlkZK6yaMaEq57KD36U5xUKlthUqP/Zrg7vq7iT9W6xeq7fmfSpQVy25z7scyy4i5PtD0
6ACIPrBEgeQmNzhGNEWXpnzYtYWQCL3DCt7RQPrsvcuaCbeD8fptU775SwR81h+ix3ZJ+fwwJvf6
W90jtPEB92XQcgJPP4tm5bhccg0K4gZmpmDT1HTVrnJ7hAAxwhhNUvOO9IiaPo+8E2L4U9GvrVtw
ELyfEbmej1f9i2V2LlQEF6+O1dUYmVaD2//Lw8icWQHa6f9OC8Q8yMNe5xxT5QW3ZB08LLHQFjGC
rQbbm8iIljcC9QQpiyAUwcV9emEu0FzKJuRxvt/da+xTOAdmBqANrtaaoqAEPzd+xHrGJu8j21++
w40Yx7FoI8UQnZ1W0SGJr9bC0xJU2Y+LWGnfhL8vTzX6tQ+x00SsWnrSiegFrQGVFMBOybgQWgjM
rM+/BD3EkbFD6p5wzDmNkBuLk5GLBXKuutQZ0OPCjw10pRLCwKlrsRoNVIydpdlYuX521FQFyUBd
IHgURBQ/K7uT7OcgsOiZEz9uXRAeBubxD0KDKxOmpcfp85OqSJI4oIEkEjDgoJcZBElbcJ4xxhIj
JX4qRfzagoWXcuKWM5pFSXCfpdymB51akKgZCRzDiE84p+3N8K9tXjBzGnVjOvcGqlWqH7Xp16tC
Jw0nC7rWIwSAmItio+RtqOHhknyhWtjfoTCIv7SyhCv2PW7y9hAVNb/GGJbA4Z+3YLvrdZfbkIe6
A/L0bJMxbTJsUaOpxm5VB3vbKdWHBZP1SYxOTjCzbXGbLGmxN5q79oBEpPJPrlMrDwpcR815wifW
pHbjPNr86lKD7bu8nAjw4IcZEhO3LzjVAPWQXNYCXZawAi2Dhni8jy3QzG4WQLW3hTwgnSlqtbY9
1Gcz3TBqdaT953TScaAbV5Ps4sf6NX0ZE0/68wby4RPJO/jzupmSOY6Quaxw3G0ic6rAOeeRhfii
dGUAg2iqS2Tp8BF++aGFwkIxdxivW2szHajK2HZ4OhU7Jf4djpy0LoAoXsVWeZQeOxg5FNyDRlvq
YUMann9XXdzfnlrvAaqQYWgBZWdg+JID/nIbdTQdJkvtNKVPwuK/4Pg0O7xM7oYTyzgO3TKTwdt3
ZvYgNE718JQFS7NdYRu3BRn9AcKufWjnVTVtzjw6W+MQyaUIIZVuF+m8BwuxEQ/Tw6syfnr+8Lbi
sRHOqCzZ6hOqFdNFXdJhzKuf6SZcVvcbqlQBJU/jK/FBHbdZT5ZzsPlznA15s23WT+1zp9yQ2jXP
PmxmH9WL3WVohGW4IJkgfW7jRj8s/56PJSvkGHfenC2iDEDOSRMwCIGhEbYuZsCW000b8GJvMLw1
og5a84qryANxiG4Bw35nJIMfiXpv+SoqFZ+STbnTTo543qfaHlwPm7DaZPbp7zRL3/56SkyP63Xo
CewygA8Sce2ur2RZPz5iP9LLbYDbmVqQqL8rN5bFvaX4t3FxndNWH4wMDh02Sl5092gu81Za+IZJ
8zMc457T90PZ0kHeXcCDvODoDus50o8cFBYtCr/RvRYlQOwk6w4APT4cAXJFb20EiSVhu6MIX4ly
7sAbD4tDqDbZ7uQm0kU/g6wOJzGWzfuwjOu8gzPXE+vZDTeMd8WGGEJeJObGSnqkGyp0IH4GuBvo
OlxCuutOlSW9pH8RaO1C8kIap/GBeeclt0bQWAhU2oWSp/p8A9/JM2XjdPg0+Wo1u7ICSA8YDdCK
qIb0OrRfXW7UX0Z2khoye/PMFpVUACPRULzuMcYOeUuT1AM54b85arG0I/viJFgPs0ROUu8vR8Iz
I4xnaL4VlXdzYdHUmSp7fw2jYfylkUk2BnDl2EcbHh+MI01I6TLVR9C3BbMWrEJsHcAhpJa7lObl
usJeqVxXjH2XqsvPK0e5RF1ZJFf0nKCBpwJ/VR7xoNVqU8rCcr3Dx7TQ6ZYEyWQObFjxZIUW/EBX
quUsl9P1AGOUCnsTfYb1ISyHykC+UlUpl/4EERmo8KAmcG4Nix/qWgeP8/vve9/i2T2/dmf49zIv
sk4t2vtnThi3Yij7GHZbGFF44oo4yJFayziAKzLIvmZK9pkdRYmMFccowEKk8gx1tudlyLdEVN4z
pKPpOvObbXm+nsQa88v6gYxkLOIV/RyjeQqELHEX0Z47uuLnxoBmwCkAmv0BRja3rGKT1JB58vZJ
4XfjrRGcP1u7XHTWx8TFrEd1ZH0T1A10SQJ0OxyydmKABLlCPjGPhBxxtU9EkunUvELsU/PpaMp2
K6uAuExIdmSkLirwdXBdiAIbxEU5MHxY6E0jQsnYQDFA5OEfW5nARG2Ov9hoTf55DaJJYqUTWfg2
LrQa0uJIKdlJSgMupvm12u+dKUexqGnLH5n3U10cQdNXAxL/tK/io7zQxvTy9lpKu8R0EqCqOnlI
f5Heephs5yKr+dgJZMsX+J3drVVhQSn0uwrrj/4krrfgaKZ9KNwJv35Mie9T+Nick5yJEvCQZ63+
ZkFY0rBTQOQOsAtj9usHTN3Ej3gl/4lPIaCH2rgta48LzyQuBTuxpYwjm5xC9Zxf42VMZXXmtsKf
kszeENnk/HlTqp6Kj5F0IJZD3UnObfh09uBfjHbCdKGftdEGDN7tZdXVkhDLesbLwk5V7x+Jk02K
eTHrIoxhx0cDHnSibvYKlH5lEaDB0rlY3QpzB/jOqHi+muObvQFDEIDP4cNB6aR1i73yzKSi9lLz
LdlBuKqYzzXGGN8LZA7NFY45wdJSrgPabySTqGSz9E65fgkzIoJl1x8nJuh5aRkIiuKFrcvFpwhi
KZI73tpMXLbKkWq7ofV/3uzB1/1epn38c8ihxTdCMPDMq/Gti1R+SEdzNxoy/szPrMeGxft64YHk
Yda1J3pDPB1oXcTkLQ2fck+3nttBLy42oeDYWLIAIxhjGZuscFVt0q/rBkaOUV290GKBhZy+gB/v
6AH+vqcqkIz7i8HgBw9EDEwj5g/gaH085SzJqjD2iWuFASD9LQEX2plm9mOzRwCIJ/ufWwNn8WOT
Tokd+k1l/r630n+kGAuSSsRQd+kbUxnOdippq0eCGBePJId312ljxoV6meestz/YaG6ZyITa5W+5
8WTz4wnVyxqneeU5CsOZ367dc8bfQ/4aQO2eK4t9X0/gyxavsP4xNaRTsYsIjBBFMy9mlJndoake
OHGHFQfY5LQIdca4UhJLtcFu7ubuWpTq5Q8QSzbY0J35yjdCxGdi6qJX51Bkcfh022LRQYXYVWaU
i0G05c6TDHrB+2CUmo9YLY/2LalcbH64aKOd492CDtWDRqqzuZAee4B5EFUWN8dG+mPgWIHhYOFy
lp4BpGxoL0eRvWZ06LmwFsBzVwCmqyIu0M9edU9vVLhtZzsZByiIGJM4ihxAkQ3hPePql3eQf/FG
U2Fk7RsueLNbbCT7zti+VNPunGA9J/DSlG67A88L1cpnDMOSwTp9ktOJPMZp7eR7l3rJPeKzLryW
1zbJncFEt1FIOv4DFjehq3bHQAsKBvkN8XotaMOnK4z9NdJZOuQugNtbLXw1rgBwgF7viIgt1hv1
u4o6KXr7nyJXdjwt2YogCdCgFoydWc6odIE3cvK/7qHYU+G4SniVqzbeUd+qti7Zyn3cLpu+lNKy
u1yLpgzNcah2QRynsACB5DprwIaydznCLUXLgD4a7qe4lln1g7S3js4bXJ+u16rQk821INJKGVmC
V3IXZdoxJTVZy2l44MrgYpbaPb1Y0FwMc+XN6Rr532TUBOX+JLyvUNSTl9LQSDIiQjG3eP7/xb/O
QuyavmixT61whLS88f2BL0kyF6m89OPxm0T4RHWff9kHVeTNFwi6dFbhUJz/WcXVlZC4UYY7/thn
bD3CQBOus2LeXYR+vZjy3rVAkc4seR6gJftSNmMjVDrFVIQal+cI6Im77svvBrSGd+t0vso4o7zi
diIBHCoHM9xY8x4qJHMXvHDwqJHdXTVk1rSMz8ih2UM2MpdJtjakNYY/O3oxYvMPg2WdMdifAa6A
5nWR5wzAV8hvVTjaWK4XY/KfW0UX1GVgR+JVape3pq5TIpGa9I/RnrvT4lU+FOJn/BG/r7dAL7Sv
u7BpU8RUxhXUoFpyg+mGSVIrugaG0Dk3oJPBmGZJ2kgCCjkQjrDR48U3KZVPy2fQa/hKXnSy4ehi
Mt3dPtTBGFpUN6BmztvNdrjGXeb97dQaKvmf7ZewiJoRXgtIB3VpGx8mDAA9+YT1rbMTSWNEaCqh
waDVQRNXE9nf87MLywxS2wS2QFSczUbNXvIj6oqsKaohrKsP9dbckiSgqG1/pBQTzV1YwL/DY8/c
0pAsO7ge78ybQowO+obqzoMKArv/3T8mAZYjrH4N4qn2+1mE+wH1q9n7/oJCaKHv8bo6CXCKPcQ9
UP/bsSQlnW/g+lCw8ZEJ+bgfqMiADxBvgumuLtbDwJPfYp+mm3lQnLryXfqpSgSTKN6LzO/jJ/Yt
zHJt6h5SVcfW4HwTbzlawTsTmboqeqV5KnnvZZcN5NRKNgZ6nQCLWJ+gjaCKWGPuzHKYzX2NZhvY
pVEDcQrBwv2aqP9j5EqG7AyEqlb1VYhMleYKDzisJMuJfyVLrHy9Y9G8a62tg2iW6ITi0tfwcXR1
u4OUWbJne21TrXMEtYQ1iEHuwKbJ4xASnzGltpc2MTObfpqOYrXos6KnXkqkDf0cp9SZUGIb4PsJ
m3EV302e4fmyv31x0Zuss/pF+8dEH0Kn/jJiwWFqLd0CwncKEs0T/vRYxUe3X7pMhLQklsnHXcpd
HXxhrS3/vonrV7o+okuaFtOm0eBUF8mbMJy2p9RHsTHcoJlSo+Pqbg7NzzXGUSWxqZnMEWtrPEoK
NIuR9J966sgRWtxJrpMCwWoo7wxVtv9E0CjqDNyt2cnyLpbyIA8xljawolIFqbZsxXO+XdXc3fxq
WXW+I4ZNiXECGFg2AIVfY18m68op4O08grykI4uOLRYY2U2nWCdHqxOSVi4bVtYyczdJAq/Hr3Mj
v+Zwpykf0hpwW7Db7SkczP4+q1XRr7V9QhveZ9K+G92TTe0wZwK3/YnPS5kq/C5I0xJvWyu8UZ5B
twWSCmXYTrXCvD0SdmBP8pDghs7FgOc0SzTPwRmssOTKLW6dPWzoeH1hzZx8AZes7td5FSaMvmdz
VHyXrx+bfvtsFP7COAutkPeYI0NDlwc541JBvUa6GXwMAtMXkf4/il8rokcT/8vRP2VDaN7PA8Q7
0uSArmN/RceTz9Y5RLtsS3CP6kmcJ4MLJjPi1NokO5bfrR4x5SfWcBeQTK8eAc9NMR5L2TIXagpz
8KSRKlxcS/hC6Bt7/FzOROq/5GkIChwco+uyzXWOOK+coq1BtrxYVqVHMfclHeMHJqFD40+8Ukvw
A0VJgXxvkBaRk0QmUE/XweLbLjOKN3L1zvUnOmDn/Pfaa/EeVW+F+jCaJlDpknUSMHXojO3QOR/0
EMt6dERntbjf4GKM8WOLxS9Xi7IZB3/ZjBbPQqsr5DjBDL+y8q0bMWZFRG3HISX0AWmb0h2A86v9
vB6d+cSSc975AOPkLKLpgJA4dWJgPPxVwNl7O9q0UD4k+9OsUiuXIU5sjDY8IAqx8od27jm+Xg43
vfNmqZbagIe1Rq1zu5hx2tz1TAQwsKdfqN/vUOVSvztSF+Kaluy1GDYM9+YcsEs0MdnPNZmsxSma
eqmzG5pgH6ITLdTVCLbfAOz6PffeZSnKfTfB0sWhehXF9jPALrultBSjczrZWBX3OrbD9yW9Y4s/
FhtVTj8vTWUqZmGOXSJd5ndH/Fb15C1Bj5S5UDyCPnLfO99MPBqPaRQTOMkHS1Od8Y0wUyd9MX7j
+UB288F1fLUyHwIG8U1vaBIOSBx7ADlcfLjMhnDMaxGl8pr6G7lw8GbGme/rQ1c5SrKbZALuAA0a
mSrBeuDxeEe2DcFroCFH7xuKVDhkjygxz+FUtFMNfdvF1tmPf5F1BMjFJ3enZd2MrrU8y34H7EGZ
16yjihN35219QyBlbxvVBEhtfgRZRF6A6c+U4lJoDNL1FtqlxjddQxYHdftx5qiB55gebSoy2aZB
XE8GRbvTckuf9OQAV8EvfeNAxRoVcpETCeLUahLAvJ+sFkjKIEaPQJQKdraG9T6DPtFOd7rybPKn
Xo2KadJ8iPBKWvXJxz0jXOYAHZ/EYUA5vcupN9R0BmY2XNY3gWeagwnNRyQOc7OY8/6F63mQEMkO
J3FQjkVJ3Laa5xjIKVXYL5ovUCf6h2zm/3mplmi9ZEg3B8luU9hLNH+RKMXc3QogYjJ2fWAasvkc
PulbkReOEUsPeU/mDLjfW3h0ZyLHFWfLp955T/8pafvJlxWkYE+bkKvn1xu3pa5BXRSUqMz0SSFI
OPh+dMfT8y5/SrkIjDgVSYf8Nzku5DJiW82doiZElHNveO1XvA4pZiVBNh/Aer5USfUXToGbUwM8
Jpqmz0kNqJ9zpERXZmcAqMy/K52F+qeqOzx0GYarfzE2b8U7GjiSo+oYgl6Yta9dXlwqxQsAz7mb
ZDF9vgrdf3gro6XtYB75J1MZpSbQkCwSh7mbrCKBqUWw0/OeLOvv5vgkiKWopraXEau+CHT0w7J/
wnrpOOGLMIIYLdz46zqi+71FBD8fHH2fbieE4LLKAa2TopG79EjVvj6ushiUaLQ9M77AzQKZdPuC
9uSC2Cl6feIo/PXJjDyfD4a9Ylxj6hvp19lBKPmJ83ohCXAYvh59MdNcmEVTMDb5WETO6b5WmqLo
K8qbkKKzFjGGGeMPuqVvGPbd3wUI7UZehsZXDy7loNGMIQOfBaudexFl8yj8InmoyEL0qezyT2YF
hVdm+pZx6V0h+6wra86Nk1BaL4rH9xCYNOEh1/UoLXGo8eDQ19JVvBONMEubQMy1i5n01XE8D5Vn
YEcIU8SyWLFYEYfUACoUDb04PBCB5bGT0Cb2+SjHWMcLjiTw4IBJu5IQnA1q19c8AO1BSrfPcH6+
HbexlEjOkRoY4sq09ObiZp1lp/m1eiu91j4jASImZJ6m6p3XjNJl0biHmF8bvOr9icu4QkmWzbcg
ECVXxudsFHQ9kYlaeST7HDXQeUDlIDf2bkbmK4CCdjpXkPK4lEthbGKYtXM7wlvRB2JmURyQsmYz
eNmZHIN0vglTSdA2V4SxvCEyzt3SFENKrO3fvBfrMatsDpGHr/tx8kJX/ybegPiWiX+KgTG8PNV6
prEISfUDkgB+J1Y9wdcg3L+dqESmCF1H1anJ8EMf09clCRL0Xtf6/jPt8pxEj2GnfDtBmrztfADC
TjxuU8LqSJBhoC+ZZgOzaePWfy2boQHVaxEchW5LKCcTmK37wq3lPeo06nEVn8O0zdY1e3Io0HRA
cyzJKy1H43M+tSiAni7nv5FcOwsJcAan73v23hh1JQhIu2JIOOU16qUlKJ5vVy+ZX1OJBgEqKZv9
Y4oTvR6hqqeB/Znfe2l0vjaRhS3VXNJNwEa7qBqrKJfB9KMAvV5ylD5K5RWZYjP83JdxmR3A+1XT
3nWPn44hOe8625ekaAGpmipqjtFBaC/C3WwVeIdhshAjCWx61u8PzIC/5JT9+Lz3v8nv3rRhBsKN
yZL26jt+naZCR4q6C0+CwWy8x4Tg6Ad/Zh8AyhwnSM5U8D2MitTqx6XxPlGVWeKlFc1UM6TzsTH4
m/sS2v89JaFBhf53Rz3p4qtt9K/+PhVeM3unSWWrht3eB0vxTffwwxXhy2Rem3Lwhq/fMhZOLPeb
9pLerpe0iLoWIuun62Ca5oYSHkGyUfloFMsH4OHzWjqqGn7u0FBqOvq+HYuwjs8uuzOSCGqxR4cI
OEUUfWGUTj3jgjLLl/68sm2GTyTDBVdX508Y0gMQDTOi7xLepepU22pCcIkUW/UpxR5yG5oJmuoy
Jy89+KMwKYPKBrUR/t1JBth3KfvOJv0j/q13w4BYfgX9KFXG6R1uWXhX6ilKfQYh6fb158iuIpM0
dQ7I7MGFAFdSk0Tk5SiA3vJ2DOW6AOp3EEzM9WGt/CXrvVnHkwhvubAW+xdQMh2HKQtKILh1+Lu2
Oh//7MicUangVyusqFWodb30admmTFaZ5pnfdg9zmqgp7/sDTgQ7UINpyOcumAb28gU6Ar26YtRB
mFjCHpwwR6C/1pPmR08FgpsnaKqfMvLv1hp1z3tK5i5utfdwtnXqydhp9xlbhsdsroVUyS9G/Gfb
zCq4olx2G+e2IulImmyN+LdWMPzXlL53/mnO34VKadKez+IVQTs1Tiz/Kw0Wol2q1CVX44v38QqM
Qb68bMaJ4DL2EdYzA/sOS3xiAzEPYsiGclJ0NWVmV2pR4vZnwgkjSEmW7ArAYXwwE2+18p2pjw0b
DX/BiXAxTsTxf2ZmxWNM6ugtkaAmGqn9I5jm/9B0qSxe7TCG+ojqcuqTA2W1bHNgobYnX1x+sGXS
yRppo6bsJ29AyfUADlsU8D244SS/Fs9kaOYy71lGLvdhYj5YUYUZQJjcTj3ShiRZaNcf5limKL2O
mE5AF9ZRmk+cJkoPLS3LzqLj1bJbcRHgld70qwx2e0dhREkq9PBU/uy7+MZWefHVmNpuwJTF8rfL
VEmdeXeCKODtG+xk2M/0nhRf/r8IMU8xC4sxWQdy8vkGVD9NvdyCmuXxK6b91pYBs+mTAsVHggc4
KRQrbSCD8rvqPnRmzj7g3xjGmgRnlafC1sYNHtEKl3aqH4ANBMMcgN2seZVx7Ua3LB//0HeGeKIt
YyoyWl7PqPCrJimYhDnt7PWzL6yj914GPNM6dhVkDD38bM98Y0XwnHsz0DGcKya2Yun1tnCYS4Cd
i25L+1a3U5hI6brUOKZDVap9GFkfKOYXZ7Sik6vjVBOALqDZaURhlOfoop88aTazRZEYALFW1O9/
Ptb1hceGD6ym06yj4APuBKazGJvIgT45b8bO9bQnl0r4LTsQCNw4GEspsEazNVB+gl+974V3subk
0WZyIunoMyKC8BEafPAB6I4A0KofOkwJTq8KwZfqifiVQGemgP6Wp8MvJRajvaUv5S0mCAVBI3vI
o3uYQgkWdngtufHzGfhDN31j8AHn/+V+103rLIsZXOFGb803n4hvQ2zj1ge+mnjbaRX42nK2Ksp6
c3qbOvpGxuJojSfdFJFSVn3IdXLtK/fFReGcUf6M863C4J0XFBkzFUCiSpGANJjrJ65ClbVZTilt
sWWhKTBAP0JEsvyLQlDZU2vlQVEa77qDNSJsd7XZj5EafgNVhObucW/SjtTfe3X4MoB1iUEnxtNt
9hSy6+eJQm49ujz65bXMvRU703E42vhtyDJIucINwkDnvaffqn4BZ02BucrAtpft4WJL+H5PfV0Z
0M2JBWMw5tl3K4jelKDsD2lpyG5X6+BiuQBTV+I/gQItivHh1EZRXmRN7EkbGkn6yQgqcgX+GlRD
1FTNecrBHb9Bmu5XEwks5o4p1+YtFDU+W2ifJxtCEc+laCbgyK+QA3wFkVg8ttM8TeJ/h9jXF84+
9+nDC17qTrx23VU3adWMgNKtoRv9q4rxY1K1s4P6R7XTUkP6IStgAYpIT0Q2H7/w5bYVAyF2Y/Mp
F6tFV/uiM99SYn8y+Wv+/3V80De9BChRG8JzoUUJMA+6SWyVMrBMCB95k2J7zjzVKJ4c/L7G55i4
dkxGJuWVV1Rev+BCeoeDI0tw/dE+XJ98iC8yGETGzZGyYiU6Dv1F/wJ7kKZNP+BHWIN1Qo2Mt6Bw
CChYzUaJcM7a0tijf9L37Xi80/pQm9k9QqzZmvl4Bb8hfdYN/MzDxnCZqT5k2v0c/I95it7I3Ybw
dzlPhOZE80T7zG7XPX5q0nIVAfn41j4EsIKaqBKWM6gFnDcBOVJBzpFwIVKMU4d/GU1OgdVzoI2a
lJqMD+L/J2lH+Qxph8B9PKxs/2q4xZvAuuAy9405aiT7MFBwRLp10eTctMIEYWg31EZ/bjcmUjeS
hESKHdnUNrhxzDVL24T9C71KmMi+UgrXrkV/LNOB5xKffAKsEjcyn+rOTt5BaIsPI993rJp4rXWL
WpbJFugnPtOnpHqBQcuDVKf9jqZ5IzJa7tCcLwHIaCg/Unhdu7dHLXmacAuHjSTvo/S3yoGJRdpG
6ssAszXO5BojsYeCu6Il4o0fZOQyjJyhNJS/BcTKT3JkoSPtnGzSH7aw7nyCfhSQCf2I5UWXBRyx
4FNzOstWK4w70IQORHaArRRZCRfkf94f2bFQVF3w0/kKgg2xQMqZJtwXsx5hMCi5Y7nrtMn924hM
TS4dJxZjnkAON+mM47Xpg6SR2pixd0NEvWwm43v7aIppQvg93Y7tEgE7UaZHxP5NqMo/qcK8ekZK
jUMBsz94+5JlLyfiuNbNKNYj+YtJ7iKa7adGSZljk2aNVmEffipzcRxRNjfkuYwYOw4yj+87f7X7
MgmV0efh2rPvz2EfvlQMwE0snGEtcsNUoz+kPQWGyvdb2M9W30GzKj0eeVkA8cII6nkSv2i7/fKN
3IYt94xe12w+8qt5zK/CKMXqyVY1OS+nKsV6/caY6nlpGWytQcssKYjzKovaamv4gay3sS5bkalt
MPMKfxPon9MFPEhVpfVf8Ye/SKKmV4LUOwWsN6TcISFAfBPDtNeCEZfkUEZ0hUkapFKHDDWVKgzr
a/mfC2yOMI7I/QlocTCt1bJMZsjtpqzgbRfOFA68iA+eebUbliQEytQg1ayMTDbO1eHAUYV7+7zM
VDG6T3P02qsvJ9BdJqJY73HmNOS2mwksdSYcmkWztJjl4ooCx0oxOcOPMygKkpwxEToQ33xhc9iB
/j2OFibJNpQAkmUVax9+LpngPi7dzKS4Fa+qNUvx5Zw43ubSE6NE6z9iL/ZZ0emSU3rkw9nLXemt
0MwbzX4oAVK3TLWdYeeA7HGiJuwcpXZ8s4lEEfopeZ6SaEZ9DPP5V4uXXGE8/nW5fQG5J9muXD7Z
qHqxqe7ypUGP/BnB5BbDRQ+J6/yzdY7fjMI/+CukJNF2QoguuTH9OrQvJT9ITQDNfrvNdR/tkWU1
7QBQjKV2a4La52KT4Jq8TFRHC6OfCV/VreKcxZyZBs5vDALEXoaH/6Qq/ULa3gUMjtUK78iGZ+x0
E09LtJ/Verh8Cr7SnVQsw6qSGoTyzHQ0bHfy9twmSpT57eCP/YYcatxNIYZgRmQwYonC+1VF5YVx
EzZl63mWP7gi7OOZaRksGpddbwE4XFX1fI0aV23riXJ01BDI1WIHSRLqprFjq4pvqjazmOQIaNbd
vyJ/NMTTgEA8vr3fw4u+fiu7G/jzfciYgw6bc5vT9ittu2mlwHKF/4o8BTxXrQKq9TJYr0tk/XF1
cjpFl3eEGlh+VFdujjPRLxm9OCiDUd5GJVrRmB8sFwj5t/hNWrUbmeTaLsJLDinWI+odVgc4KLBM
YXSATQW/euGcvvIcFroH2oQW2et4XMiP05bKtFAe9JphZTVzGEM5UjP4RQcRlgKhpEMmAHoF6tcr
6eslkWaD+FKV/RMWITYREvx7rys9nohJijKSF2RCQUUu5UBQ57SVjTMZ1RF2pONVneTp+D6j+Zi7
s84B4OMK14zoQbKWkGR2AmqCQUNDEsH1EpFs9bGa8ixfutNcIUGS8U1/5TWA6Ye3j0+jZaBRSUOf
i+wVCyrNB2n6swex7ClLi9yqhYlAo3B8GxZPJJ1TBEQ0Fw1Hb29e4XIJZRGN1PALF5BwAwCbMx5f
nPn/uqc4AHtGWjhBlz0GSGwRcbHXEabrrzERVYScOJ1Uh108o1rToACHDKx9fJtLGs9bxGeWoYb6
g6b+nS0XIEpXVotHUsS1aXlFn/qalgekus0no4femkZBWWklfIi5OiesoesUFXwEn7KuDfKEYPO/
Z6AeHzPubdlMDKdGFgOEFasA9WNFjghjhbh6tiEFQP8Kh+H4mU9bUGia4uisxplkmXym6AuA/Elz
kjnghHSb5zZL38fxN8mXzGvL/yKYC1JH4KWlnnLSV25LcW4Csr8hjTQsP9Z3HNCgXIFl/95rDBbp
rQyX6On2cVgMdycgsKQRsnHyCXn5YOqciJ+xyRUnPagwNtmaQDz7cTaC31fV1hMW/H/VuSE0Np8b
OOGJe/qo7o8dCc/GomqIHVhYNiFXQgYiJKpyUTryescMv2SBS8ePal+AYX87QJj0QwiF13cEfYIT
lAcNWeaJO8WanZM2VLzhX0sM1rsQInH3hQXw+0VIIUnDdvMEBTv9YO83BCOoCf5g3TDjTcSDk1DV
MqPSWxO1ePelq3pT0n3dKZxzqUhifEZbimJPDfRwbKd/8LP8mM2uWY1rO84nJMNg7i6GH1jQZs6T
EYrywYx1ZCUbQvnmS09SNpmwG/sdn61F+csBCR8Q04xKOoe/DgNpCrTusxTsfKSUU4CoQJSBp3OV
lCJOcUVCcfwb1fy1aZI8o+IcoFIbya1TJGhOjLA8ggo/PZy49ZCnapK8eJJaz1oomGFrqITl/QhB
vl1qbJ35ztuWRT0OqW/PGPWl7cebaKMQdtmV0+uZHn5+QLJ5SJrt8BkVxm3T9E8aw0d3hySYbRQ5
MGai/e8eFQeyNC62GrOkHDHV6MsrJJ+vBenNGrz1tSxc5611NOocyzBhrGpjJ/k2qraZ1qKHWka3
6CngGd5ag2CdFXppCs1NX8cE4FTOkoRpzm+iabXjWzuiYgBFPb/4+5LTTMSM3DYiwbD4dVoVWlSF
RYMAHX/Z0/jpGzSCOAsnwsritv3kvpgxGFdhJHzVCN1wjAQss0FEthOF2WdH24n8ALbsnGv1xGbE
sbbhzl8KbaKtRJtvQeoHcBSg/IyV3cJArkNKzLhwG4BhwnVAJAv82UNVt1kNYt9mSYu3OGHK9ZbU
PDYkARrwIntpq4QVml9R2Jjw9mgogHwgoBA9l8AnZD5j5DKcwRpAfhVtpTG1kbBcu8BQZxxxRPs5
zPlrFYs7sXAtTGm2bJBIJnkcPr1psF0RZeCx3J3DIQuKJ63F6zD+Nlgr5fIDEScXMKWP4+F4ZAv4
RK0zXaLRiDdU/wAoTXXKuAWeyqPmllIN+UfQJ4mO/er0PpXCuLOi5At5KvIIiPVbz9n5YGzV81IQ
9eyv+8emA55R2gNb0aF3hpGerQMnvh0pm1F9izZ5YmL6vzqsJ/G143+fh3PiqqMcptm3FQRYEn90
CXMLm7yzaXMpEwB4nIwMNWu3t8aGnkNf7suWk81jI+qyVA9ciHr6pDr3kDjeEhzheSoV7bpgbgwh
yVZL/nSOKBFpJSyGGkCOY9/L/hfMeBV3890TTIfWAj8sqpXRokPqG0xjdZWs0ur3/WGQBDOkPD35
qMvP59Bxn2oDZdJnhj6FA8BDhxjqwJDjYtjb5nMsUDxZyccYyZUReq9tDZoSVQCBs5JIAE7AgsVg
Jo9Oscwib4oQJUxTon3/bUgAChcPhdR4krPARaZF1Yko+s+I+RCrESSjQNw18TL/kTZwzaEq4s69
v4PyOFZHwTzkV7PNxXOeQb0yjT7lZr/Le4SFDWItMc70BMNNst6BjqCEFtTHTmLe3m+/soR177Hp
zwGdUl3VhLPbIyskhV+yZ3a8FG4cjRrVT09IWCLn4RIo1BkgDGcnNpk8HDvtMZDdfhKSyNeDCu+U
rRToELj/xMevSBu0Hh17ommhpnZDhRvi0ggebpxqLSZ1J5sKcjPVmmrhHIBe8GPiUG8G7hnMYIqC
qBii8d1kvwNWufYS+Wt0BWZLqQn77BFqidDsrhagUkqPousoaUXrbzeQdXqzUwqqGRKtOSF47gpK
R1tBZuV9FvzP59IJLAieVSnLW2uINfoeAcVK0NycnwngvKLpHskCQiXNRUVjXINsSQqeXa+GZmxI
nELt5XCm3Q/Tq2wSSwa7cKMxOP3z4b/HVi+ajBsv8WeZx4jbLZrim2QUJNWHr09tW1Z8443AFB2T
mgUMsc9QIKiOi33fi6X5DFDRFvSRzASDd/1H/iErRfQ707KPvcvp/ElYkjyJXlaK75BsroyvipIR
O9nIJmVFWwjw4RFrq9fS0esaf1wRwcwQr3s9vE5HQQk4CPJuOEhBuuuVxWKfHA2RyCtrYflbb1Jh
FtOsgKohj73J20goPwL7R0b+oRa+DanCcV7M6oaKVn/qBn8UIfjLxmwrayLy3OVuF8zsrOPJlOIk
hVYua204LpQqtwWSb0yovd4I6HRTX1/aQqwKEsddhBFOp9fl+FWk9sg4lk5GFNj7WR0m4VxLhSQS
JD12yl6PUffxVnGWT2jbmy5eAH864MWfJ7AGNf/yODGV2irTDSoIz/gLMzu9qFgWAl6ha4isOk8m
57zGqh0qt7XS7CA2TQ/+kjXX1LdAznY1oEGTny1PtZ7AMkUgvsGRYd41SbMEVS10z4yub/jJX7Kq
UoZAc1a9VzFtoN/sSJFDtqHA5wz+G7vF8vymLWHcKCN6bZ/8gxhg1sGZahga1sr4Sk9YxeupQt2T
Iqo0fpMj7sr9KDwudKRmUTPog+W2Hkj3AZi5Ow0877Vl4j1RtO0ULhPKQO5BjZ9Pum6t5el4c4FM
xWTyVtkc6b1FCeY3n65zWbPn4mbSaVbjRaOu7gwzWxlbBHuzjm2sHvrDEdhGZr4XTNg/sKzT/Y5T
wR2kHz76v+Xh+ZoABuQSS2GHTEft7eMrTPqy187Dwc2O9RNsFKrrj6vOFSFSNMsn5h+ZXv7QyqJq
2jXIVly/attdvTTA4MNRM1UX00iWi2XGJ1XNCgcZmTD6ch6MjGA5azm38bVKN+6cJYrFPkdv7gYB
Jnu9nwtciQj4AqW+afh7quvjHmyzF4NVC9iCwkMSC0an3EjiSDukmcvEovLfofZYVYsWgX/Q5XI+
XwOXkG9ldmLZzRQMRv5nUt50lEg5LKMhbn+dr/x7Z2fKAFmvwjCaOt6rkaNqH4HqJsIMRp15tM0d
7aXOcSagalRYb98R4vj4CHEQoRyAtT8xKSiOVlH8zo7bn2UE6lmHmruxmjC63eIxScX/pP6c05ub
/pupPxa566QA/HTQiC33QIN7esVqMhXngIsaxXDba1PF2cwUbJP3C8vNhlnJxat+dVy0qxD16i2y
2/z0Do8paGje05/V4PYKyyLW6mfmjPCPTiX7csSUFicPFw2oZ/rfqfqkiDpjPMRcubNpc9Gp/jL7
QSF4H+bcLic+ViEPRyntY19Iriyxq6nXApkgjq1Xfhijqc1Ff9TZVcjyQbwAwH+U6z3eRBo9x9QD
/vKhdtPmry+TUVQXSdLKHXiFQM381Kthotk5A60qH8xfDmYMkWNOBXcCGQ8vZeJtVsYroqk+z5V+
T3HIFobWwci+05kWlrCB28i/4vCSEbffplmUEApHTmCPixOckZDqoJnYwjgE0PEgaZDx60SAsTz2
APYP7cen7Av9TV9aPxqDWhELelo9Y/QLpJqBTYzA9CjPSJ/DIKgiwaje3TDN1qSQqu/ju4KX6u/k
+ItEJWHiZLdDGrOLwdVDyxJm1OdDIppp+K7iJKWaV1CCN5VFCIWskhZdRbGip5hsT8DBwb6TrDXO
cRt7cjVky7WDdrens3vqz1xcjywu8j/h9vmOFTYTBeDosAWeVq5YLQxR/Z7XgmSJg/10eSOqyWBF
yCXvaa06HMeUCTTkBtmNHsDFwnT+To7N3k2sI3C5vXdqGUUXuddDN39NCttyiPWp5+7iOvZsK1Fc
637yXc+yX4O5PWZ7oHMqowTdv2DRnh9H9zsmfret3pJPojWhfCBCwz7h9psTnSEWxInIrkxpraYg
Kcuxbcw4itOHq+9x846ATBSFlNxoROyxmQ7VH280UgOIeU9zSwSAqfbm+rwsmd8zzMcJh8iK5izI
6hqSSm/dPY2su8RhCVbyWlSx+xVWZUbW7khSjZmrhggJJM98F0cB949wxTCndJp63iCgYDjvKmQ8
dCEE6msNLc8BKBDuLz3Ajiu/4X4P6Yuy7OA9lMZai5PyC2f9kce36bdT8XVKhx1hSUpVpT17PbSg
39WSs3AgbrYPnd2jM4rWPiyS8MfaaKq8OoHuQNbkEP/sgcyzgN3wHeV9tMlaaaJKWKWF8AyfwVlN
vENFu5I1NBL07/OZFL8YJOpS73SN9Q8AO/ES6wjKAUeoSuxPkvHVhvEIRzuMEvrOpWMniqCq+vaw
RcwDDnDpRMuRXv6N9ArYtn2K2HzTx+CpXO4FQ2CvSzMdsz/FfCjuC6Lfjaz6eHxMuD8zb0escDt5
aiw7V2p3yg26Gx3idMpWe+QoUu79Nt3g0TxNfKLB4vA72RzsJPF3yFGfvit2TXJL+hurLXzWHaVd
9QTNh5ZjKtiWmJzAXmZ9UrtEaGazcTJFOkgMzWVcx9VwN1OXjYl156tmiccCi/Ns4sWvrMigXINs
JUY6LMDFK1eFsvc7C4fMADGqvfrNaIb/66mabW2yyWSRTPtTls425fe48c/jhnyEGfYXEN7HSDGk
T/MeSIooBgaTIlftgacGsGZT96/GKDe9DWfscRwMD2r2cdEuMtNHxADuhicGXNGNneTLEBQwOPwD
GmICujstQL5Sm6af2UWxmInMQTV9iVKv1saQ9nmQQqKa4dwXDJfzy07rMvBMf3qvQm7p9XPVqJCS
RevlHjWvxjmEYxbzZLkVt6NDXUI2dpzG6O6DAAVG2d4w+UYjtTpYMGzaPh6EhHIq2foMhrD7rKvI
1AgxzSfrw/vkEHsXvzt8k56DWju0AUS8hPyGyArldIMSvZvKj/nEv6tnxE4eJRc4JCmBDh8nYlTQ
pUQnpUvC/rvKxSztbSg7H/jyC3hTlBnQmyZ57657Bi38WJYt7HeJdvbOn6NccjNiVaLnh6+VVEU3
emKfr+k6zmRJIZIgdPIbhf98gHhiVdM2PjRbyZujZFFev4KEPqbEqZ3dhHm5LeI3/KT9sfj7QpIc
3C+6UDDEC55h/GH+K7CtAeaBiYiadH8rX2Mai1Evr/ezFCqf4sIpbZsIZKK1wnLOQeSpjGvbme3C
P1dKoXxgpT+0y489y+EhKyTRASEMGNMjh4iu3NRcL6rrmfNnQSZzTPZBj36NWg8rDsi4AmhfJH4I
A7t17z73PmV/urjY4xEckt9qvXtolgMQt6qFbtGoc3nYJBRhEBH01gqVeoUTAdN6ceR8UOAd+Au/
f97nTL6Zc8tRs5vXtgFDlhZ3IkbzBn2tVg15gBYQfwogtyRL4T0sZmTpqkNUldc2immXEfYGLYdh
QPqdXuSL2mHlj9FqvHrJ+98Rfe4ssF1gKiCGJjUb1pNDQK9SBbIZ2XoyD8wqLdCZDgEBf6HVCc4P
syWw8+ZqwSjUX/OJ5y95OfVAhk0fdcvQlGakjsDc2oXbqRrOlAOUc3pcBuNwhKWXIBkXTkrhzVeT
nDHXt431j1TWaDrALhy4HeKpe4r3pyGkQBg1YjDwL1M98dVPDNTyTRxJnm9SoeDzoSMeWaKTSsu9
nKU5388ktrHZk9xZBFvRj0fjCGFSFfRDTDSsqmsnBbqVK2ZFnLcrl/4Zr8VHEi/7auo0YI5lC042
pQLUIvqOYxDtJrKuNwNwklV3HJtOZoptbzaTVdPGBuG9jqgNRyryA3acuqf+fYIkMgz1wSkNo339
3Z6X1OJu53gK0hD2HNrf2T/sNxtSiWUGn6PHviwUO2Vj/8IPLwgN0FgEYsBfQkdAdtEsDvauqXue
o0bgYyKdugnIigjZhon0I7fZauy2LhaMsAOJkP7og9kUnp1YOu/t0QGMonN/9Q/4RJB9iNggQaDI
gjladNx7fqqI3vpCOKvw6ndkmKLxzNXACUz0SdQpmcAL9O6m62DhDK0gxvOmNVXjuyUEyoeEMAFf
P1MwJMC9fixKtbRxAKE6s/8JJNOm8u6s8C7MT5Ed+Ky/IrHsR6cmil8e2Mb2qnIj10cU06b/h0yY
2ipooWVN8OMVqwIlsoBM8ugSQpiAl+uP4q05Eae+LNe8Hqvcv9aH0apYncS7RQb6DGJ9aWKQ00lj
wCAsUr8cs+yTBByutEpGprWQGvAfFzuNN5d3Tet0ARkzIVzhNcYLkgvK/yCThQ3hP7Y1+4wTLE2b
3AP6vJoahjDjlxAejdCwiJYi4DB5FUtt5uC3+VZQTW5vqUynx7dlbPSa9DtbGtbkmU++cdOTOCM8
BQgttsBOvi/NVtGNu5jOuiD+hOG7sNTw8pCoO/b8M87iiuiFiWMmzTsBuEdyaIwmdZ2GkbP5yd+o
KTXxUeiFLRbtvToqv37OiqjAMI87Y5wlyS8hBdrRppFvxK36V0Vj/SB1fIoyl21HOhNuVqf9wmVH
GfZUo+QIQkWCobmE+cnsUrOvVuZbQqato7HvVNZ3eHIOmcqfpveh//D1vjrugey5PYIkpbG8gmTg
7JxyTbnUneLdVYYBhpMs+VP/XheLzKL33hNNr7sI7EH0M6qlHKof49azih+IVRSwSQcgBgBKBUd8
fSSCKKARz7fgEfJEJV0c87/URbrccC4bOxSbmUxuOqoTFW5Ld09WxZEVVHiyVd1Hqo43rJT353tt
eSIuJkBftJ3Fo/DTb2mMPuURhbpyme3uH584y5l9k5U6xRwgnJ+UdrV7+PDb9baPxFwhoLIFrSl6
uAgWMzCxtv2MDuNdGDBTRaaX2v6tOsO5SCtr3lG7m6JfM8MzFrN7kS7DYRXA2G3bbwIlMDk+325Q
rz/A2uyPmXCrTADf42Gf55Bk5AG2/Ym3l//SmU8Xto/jD1xEj16D9xCHstH/gsTXcJmiS3mHXlg/
2cSqHH93u68qS0vf4Vl/qyrWJO1tuZ2ezX/Pr1VdgsOanIFNk6gbsg8isDN0tpG3nOODMPibs4Jn
VUF6wzpAW/KCy3n9SUItr1U0haVc69DsVFrztuOouyzUkzmELfvvF5iJirebyD/TV3iSqZ1XIO0B
I+iEi4JNNc6BUZN+nS8bz0TksIuYrUHYDS1CWK/X54KmYpn7lY0dhIE5Y5ES9jsac07PaUBC4rZM
4Eg8aSJ+8wWEhJsQhyzWu1ostfO+WydehEL19WeQOlrKD/2EervIxECCdOSu2OHRkcciAv1mNDzR
7s4Jlxh1wKm6HeN1DSyR9rRJGIx3z8SZoFUH9yQgE3gTEkPGfU9m7IE5fMm+i2M6BckPqAY0yMQ6
FfjWdOsHBm6u7apdFzQ5g9ieV1Jk4eT0RATT49My+87/16QxUpCUm4f6trgpWKrfjp/lYk26VOUm
foonqb/Qmh4mBTxvRzOP9bgEaA8sAo8frs4Aij5CIbRVyse5XZapZvuYU1iUxUXP5lSVJmO5H/+C
jOeLBu0y2y8geHtn5j/D2jPmO1RO29fa2HKd6q8hfWXddFjQO6Y67+Q+ypXaIC6saOT513vdEckj
oCPhzbLBG6qRqLY6JdIp75FVME8K3tevoejW1rGTea2ElgZER5M2JJEWVFg+H6U893GGlCzS+4fu
uzpoQFbDn9yrMWQ5kf1wDYdZ0vqGuIfHCYPAXhVSUU/OXfl4GGsuV+GzIcL/L+3IGJBX+fNY7B5S
30ltk3o8iVwIgDygZWK6rtrJ0rK89Us5sNDNKrK0sHIS8j10nPywRdyDSQh3IUWkBb3ALTJ3MeMj
UYhyiUMFAw4rfVzNlGtIhDL+J6rtLvsxuZX79WG66iovO1v9Yu/nNVVK53fd4/uKyUOVZFnz1YUo
0TO9BvBWieskxPYvTOu0gFXbIrtyVEwDFNLpPKgseSeDPofJLJgc3iF1ZDlt/DJLxSSTsifwSpAs
QJ3EJL/D3+EzpQnxNxif3JbG9/E5p++V1v2w41GhB9nhdKHTt1ff+IxJ2ZDUXBnlNGrqClJUnzs+
WX/lA6bnkS6uDub4jIwc2zH+SrQM5KX+UPbS0j6Fnx+OWexpe6XzrkTvRCRnuaC+P8eMdQTZ79gA
+itQK+IrxtxMXGHdWDPbriYEQAgqXVZKdRXIask5xedDgUYQvPnjkHZXTB+9KImYLlCdDG0RQ/O2
MB3hGDG1XEvG783od9TWSBq5ztvTlxJo8BpoQ7lWypIBwe1u5e7RJkav2bneY5di01ugQtRAMSym
WkJqyTFeKhmHMGKH19oqzdz5kpRWhg+c7reLBypmjAAMdFMsccm788noR20PBjjwhWzhAenHJm6d
s5xXF6JtpyP0tsVd9u5Esk2Rbav9FyDQR0oob8cIa9GOlsTUfyiQSCh7vWbCBBMbU/YJAbidVenS
YcUnOvQ7rTgXy/sFctnSHqXuglvv2Jt6LvliVmr1GLrdebttmrW6yV7zRCX8r7qgSv/IMEQt4egy
2UjAecuXoTPca/kZVT2m0+Ao3+kT4DzUAbTvt/JLqac5JDAWtFq80R8VKCa8f/XA0f8DAVvERgon
GUOwMZEcnnpvyrYaKEknm4Y2lncatAQAxUQzXlewZAiPY305a9NwWXgNSRDSejL1jYx+bO8Dn6Sw
qCozd/zVe8cq1HZBXDZZ+7RwALdd5/7rds44uI7ZDQIZDtn1Hh9twYr6nsdR0qDzUa3vzcDfJP1E
izA+ZLjYouaLTBs7T7mzAVLOozbdGutSOX4drGWHp1DkioIPY9NshyNB+2FDK/QFDbogc954Pukd
ojXzkC7soZrHsn2pF6Zwn8IO2puHRohGpXMvYmZGBZxSmgGaNBjl7IvXElP5dWAJDsz5dALgQGgv
LKMWDUuCZBgYzpE4QAs6ER97BzQF4RCLbmcQ4vciYLBfl5p3cAbzaf6eW8lDVaD5TQ7BSBbGPFQK
hAWGLFV77DkCFEKeCQh3Ev5eM8ZG83SpfnJ0iGmc7+S+Zokdiv1LBS4xP82LQkc6KQysEs+K0Zh2
sD9Xn8OBa7Xqxm56C1fRcT7snX6vpXX9u7uZh+ZIHesS0gXiXQm8ZLQSuRBnZsdty9Q2qBtp+xLO
9FL7AG8B2tHmtHA6FVDfi2RTL9Pnewc3Fv79I1EBi6b423WBKqa9VHTzUurboYgTgXQtEG/M2aDC
NXiQr64sOL3bWEkjlHfDtFKCVIUIYDyjXzFf+KqE9MReNX70sEwMXfAlSm6RLs4ljk4ZVQ6nLsvl
kxDnMjHqUPOK05XSFOJOWX4WlS9udEwI0m8wHGTw3+sGqhIpCjKso3wSkSV79hNWBKlEB7ZRpVtt
pB4rH3Sd8TLF2nmNXL+uqdys1wn8uNsQqiO+nka89T2umaDzjzQjV34bropBQuwCsurq5KlFeCQ+
VBtLVXzV/cc6Bcp8kt+0Vq3VKw6W0ToCquHSOX4oEGJ1wr11xXvMm9dtDqOwhMsM8rYB2xutxxUE
63yzkAy4ueSNa6NdbOKApOhlL3KWRh3OWsE6WglCt3W1mzDABF4uztR4/QjkDWnHrFnlUyJHVtPD
46FgR76ka/Sl23AI3Gt2iSN2K86stQw8O5Mh6fZVknbDapuFQocLMqxhHJdxtUe6GOx9MjSuAjG/
xuuhBvyMrqLCQNiMsLZGe6TVL9lnhh8Gw0AWOSnlWImanP8uX1YqItI3lbTlXfa2PxDMZ7VdYG4q
/bddDboYedMz6SHSu18eK7gBrBNsPt3WnFt9Y2tVZhlj5jy09KxUFsYxYItnvfHO0nDCGGBG31ap
EGTn0qxS2YCxWo53Y8+LnzVVuimtJbDbRvQdJzuGTnWcQWuIeGzOXg1B+CivDqeB655Ah1ewClHD
IP0x8TMl1tyVDxeNlUeOW0dN7wf1/3m8Jq/QWDdz3XbZsyZO502Ablz5XHYgErcsWqEoZEyHziOA
lJttXLMnYqoQ287wzc4VfrALPngNIgUBHgbPwne/R2TN+s2ksxlTBOU+yeXHOYHR/3+ngPoc1g6w
EG0MRzTdvTPA0RMaNQj+fvYcZ+M3HxB1HsBp6Btw45VekuJ4QKgXoqOhclGgCyhmP8sw155Ul3Sy
M5lJ+urWGSkMKgr5YO05+A4XSM4R3Lv1wgC89ORVeLGulDdqeusKbpocLg9rnXDEcSX6g/RFYqer
g6Ngjdu9va3GK4qI1QejIqqQUxsQW3Ksn8XK8nfye9bMO5xNTxjmslTHgHBC3R7ugx30EnP0ER2M
sGYUhW5XiLIkDg0EPR5SoYFcJpG2hnt20salMEf6bKS2TyeZSWwU1LAqE0uH5v+Yc5j/GQ1B6JVO
pzZuErSPT+OKKt2YXpAEA5jZTAo+QA3cYeyRsFmkcPd4P8WAa4q3IB9PiOgtVuR9taH/s7Zzbym3
xLnEgJPVcSkjvOdTyeV7YUAu9swKVJS24CFGzf7x+t57f4HjOTu6IqZk8nl33vzTFEHDR6cfRPsR
TMRBxI72Q4Ib4BC0kyChwjS6ToELPC7jqVPOgpZEOmpXFoIAsIUlj5dEk9UaE7rvy87zJOjDFOeG
GaqmV+guXpkoWrdq3DELns7QLtyLLxXBt1z+hVkW5Fn9zNVqqigC+VW9PcZnzpMduKbm50lBHMOc
II7fiEHNzcwU8Ee/Nbqoxef+FMt4BFG8LaaRFMCyKivE4QNGOShNyEWvmiDOT9UIc1NLScuzcqVL
Crg58wrH6QR2YxlUGFxnIx9iK3Vhzk3kqPwjDNy699QruuR6ThpX8jKQXSBfusWqO2VLrBytEuHY
iOzZaWo5c5nykMCjkBRt6wGELTXHoOymxUaxBp0LLGmyjJZgvZzeNAtTOJWVkUqq9W5b3gZo7ff1
TaIxb10Io+3bXWwpHHGhFsVGRAthfjDtYWhFlb8WTENKLYp/bRRj9D5ebDnQmfKM81vjbEGYlpr+
Z2eBbHDKv46QgqnOvMLurnsfocFWKgVuoZTXY68Lw+nCG4ZWEB5qQ5w2Wjyrlk8kYORxfl2eLwsy
aKNU78nEqmdfnWIkd+rMViLtcAcv6fDHTx6h5d2XmAOG838K7sF078dp/+BzYSfPrMe0zc6WucpD
2HSTaSN41b/UJnlNa5b3UqyImmv0VfBFFkfyTtCGN/So0BytIuNMkWhm9SX4K6KQH0m2WzIrwYft
NNPM4LJE+WE+HcxUc6C53ZuoEPcKP1tqnjzulVzQrBTcxoMdKmQNZq10zB2Xyy2PeDg58mZL/HbV
AHVKfRUxSDEYA8KqLzEl9gRjSJbV8T8Hvuz8zCe7XjCqYq4uTzgOKRYkmlvjQBNSZGfBSDq0yGws
gMMvrA+SOKTuQtIWA8uqzc8iAWo7Hhq+5jdGcBN/7AoXrKCDoT7X4SB+bpUdrQpQvlPae+8J3GKi
c9hoqSh1QYjWByNJmr3wYwp+MzgPNHtK8DOFHRs5c+UakNMBiRMGT6J3PRdHU/RwtOsDNtIWmPiu
a3ZK3fSzirwes9hzBvBAU4P7FYWrk/DAP08VHlVRIdmo7x9W2zOK0/fPRUg8aAROaMZdGX/PYfMk
rCO7TtK4cGXV/GxhRYGDBkfS38rOwcV7Me5pRgFABdHMAby8JzdVhXipFniFiB4bZb/vaU3yDmuw
yNoqZk+3tyJd+/gOOJ+9+QBvCZwx71SXMZlcPmTl8p/ioDYKV5MqWLjyN36mxYWnXgwh0TgUMBwc
QnvrmgHOrlxXiGL60fhsL6k+G2XPLGeW1q2pon3FjrrcXfcW/DIyZV9ZGL4GY98nki/e2+74PKdE
Wvp+dLh3SMtVFMIjRnJw8oX5fQcwkOo8rWOvnLUCzSv09qyMrfO6O+SFvLGnXS/lHCd9AZeD1uyP
6MpZOYeLwFuT7phLxQ7bfz7BEQ6k38UCfljpzxigGlfvNXUx4bCklgGDOAEJp86d3DNAaPAGCu39
UAUIybFhy3pRNq04mUMjwJYbseaJXRVCz9youYktlFbLEUKpLyuO/P2NanyBJuGtpx732LGhi+Ux
Nx4naXDPrxwF+ZKvn0FLnLcohg4yNTwyMc346x5n+rbyznm+n+vNfIvgkYSo+urPqcJ/A8lEBPDJ
4Z0CjQ1XGVRVymeszRheY+EZtvzj13bar3BigqKety4MuvIGnFH1JeLG+ORaB6zPdx5KE8XLddXs
lvlOGkq0xwkPsAiD7FZHAE1E8JQlna4xJqH+ai4wFER3C1NB6/z6/5L48B5qeKLpR9BidPzZsbnM
JrqC3sJIW8taAXRRsRsNHHFjp5XpvSLarP3p1ugc7gEztqWSYGlSGv+N5WRY6xwxcoxG5uPDWBQx
LI1ZUjg6VPRlabV9CH9mTYyTYJXhCJxbxwjfZP+YRZTLuPHOqwT1T8A6BWYOS4Te6ykFTHfLP4lu
mHEOFAPmbNgC9jwxU/vuJeotbBnEz7JwHZhinYLnbpHP1nbuhVbf35CIiAdOcRiPRJbI4XbadAcv
LcL0vlXeP6h+Bbrqf9fPgMeUwi9LXkZR/twrdPDgY4NGYVJUnh1BR9bguUTxgOjiw1RBNMnwIcGj
WYmNn3xPWMhmAMi2zhKCVJa/EqAbt9BJMMmJMQnxzGmQd0ySNcB9+cz5uF2lb9ldJn8AL+ftv6/r
ciIw7WAIXSfGdKVuNL3kyOPgc68I5TW2vkWtGOKfa3Kz6Yhw0+y0dT61eRD7rfP7IrRNv0DONAFF
Ydcdhxjo0knssI6oNBKOx7nJ0ptGC3N529Bl4sbJA7vKW0MTPuuFfybBWoWav2osquB+Uq1tOAwb
gX2CYzmNzEszlItpzc5j6N+tHs3r9h7+4CWSobLHPfaKXXiWzh9zqs3ud3YgBGTrnIAaXA0I6Kga
77lr39VzRN+ItXMI16kQO9VsldCCIrP2mPEKezD8SMgyC/UtK4BdQ7lToYAdUBIowljofQPwgzIx
eMM8xz+i4PkFzjWawMVONe2Ue33+rTESUqCTxOjrBCpPtf+o3CoN185I2gOEbtU9rpZ2CA4CnhgC
5IemPJxSBBxwbd5kni7uTeZKZoKpRRdaoMYzK49gpKAvAKeS61wzf2XsSAy6dDmsds/cocfFeYok
TIURQxIjRcW4Rc4hgO2VPHk+8lMImDqDjex6mels/rmK05YMJA7KZ4IWLCphHdgRQpKPMyO3TfJR
gU6csGFfXjL9csBKazKHdeNOlLqRGdslYVffLf0Yx+nkVeLs7LQz/f6NM3xmJAioxmmbiFzmXBin
JZ4jCQHezBMgKWjxTqndtBTkn+P3sm8ZrmPYxvYDSracih+I+gFOXEjirHbfqhHHbYYFAfGmApdr
vdZAPBcjuXqCF49XmSfEKJcR7jNdFJgXC1MlPOj5aaYic2d/tkjor4zv5LY0OITGtf/R7S6aLiX1
IXmMA1v3NixUq2R7P7UN+hu3v1D3/nok8Y348XA8gaRC0mFds/V69cWHdGrznCbJUy97EnRb1EkS
e5VXwv1F/OfN6rgVhu0ce6NjvaBNOOXgcYfyIkTpAm/TfYX4CSdns02cwsweol7f2wCMuTA4M1oW
cR2WTeOl3bfJjAPWGmsBJcso4OyONuxv4S5IIYDLli3PYNmMRO6qmo9XU7r1GHO4F0sUOfFPxS9l
JRg3NL3EgMNKbYX0wv6PLGOzbdLd2IYbRghRuEcpuhH/S8dCj9UFezct/GmLJRFQHdBCqY+4THD4
b29Nr2tZlLjTiYmFcU7QxJEaeXsa73dZbzWtcI68GSYzb9ur5OBIlVJ5gAosyCfnkVmhH5FZNtiY
3fUYlCLqjqcthE/h8hZHTV9Uq7IlznwTZBEqUrn0jhQq/TYAcEEtfTbxE9CEOpxu/c64VZ6X8BKf
fAQphJhWuBzYD/mzsrlbRm/tS5g/U894M61htLMNlmMGM4oG8kQ5xt945XROeX3ZhOMsFin1ApDo
8FObQBwNNXDdpRtlVh4MQ+5TgdAYKNXZPBhL9aXTaMK8kYl6gpzd2/Qci91pPGW8MdXtxUl6Zy/d
B3QSXGwhAU0ipAl4uynDeKkPpwFGeIvZSFRTsPOmNiRBJsTUWw592St9OjyQhgneBw1QBHjyyXal
0mleO9jLX47D+woMWvSyK3F+FB5UiQ7W6X2jUs+w4FeoKSYpW0MgkwwXXVQ9vyUf6Di9syzlA23d
gIrLdyUIHigS3wMYJq5X1wX4L5jkrxHsUP9KJmV2Zgb5cyTPiwCNjM9L/1wnWUiU//5ALAdzRFzv
NGflf6hb6X9bfYlZnOO8HpQNk5EHGxXIFsxh2QljNjwPsRuyjnt8Ts5tAiKgkTIc9G6tBRAg43d9
pjuVcmKiHekk05IhmA2z+8vOfe6NfJ6JsoRqvPKeTpJo4A6A5VCbEBJB2O7aMneuJHOy4Sd/Y1ei
U1D1vtuOTpY1n73F+KIRrvsVHnNCRRvNPoM3GdzXhUvYB9J6O/dBcSMjbn0tJt+RvlX7ijvMKzbW
KhrF/mIYWq5VCtwHrhFDZqUrPGaa58NbWBG2e6HbL0rwMKp5cA0wDNc/oNXk8jh7McLQNYG0TOXq
qBnoLDrqbdrfoXdUWWFpSZSQktZ1goDHzI7D53PGv+2QJ7Bx62zWgPvuotf1KaJnlXwypnYPJFS2
FoalEEPZIzWTyOejYnvNF9KL0jlj0fAr5DNh2muXPmbAIgmcTKcJcqv5rt7C5jPCx+nfPE/kW+t+
IvKD7Hlt3RExm36aIuWhhyfcEgpIGyhNmwh10NicXJhlU00FdryHS7PtyZXUf7AwpOfW9ulbr5m1
n9nKnZs6EJOpegLWbBlSm33wOKcfl5e0M5LpnCSvxdLLbEo8/rWCG6ys5VabSozyCv2QfBT9/NQF
fcxvSrJ9aoWovTC5QvsrDvN9iJwClepaS6wwxn1yNSWzW8NT8xBF9NgoitxLFc3mUsHMHqTlXyqe
/zpTZfKvPIAphy0R//Yn+NT7ZeZ/fODDJiTkLNU9V5y9sjnT0Yl9EqXW/WENCWJyT2XdAgcaNnPj
RtZwQX1rWxEY+2iePemVn2n3V2GJJ6IZ6PliFKDh6iRyJaH58HmaZGpHP0bzoUyT0To55R7jxgLg
C9uYEEyq6JwDOXfkUK2g6nFEi1a2qUj/qXnfJAcYM50A2FfpYZIcQ2uyGe/qOckkprg3PbzQdcsX
zHes4EG4fN/Y5md65C+IiIfeHFEouqtMUcRa84qN27VDLeGWzbuAPXIALeVTeV7+0h8zsUE8I51Q
ChX3aMUe7L1zCK/tpi6J+exi7sE5Sg1YBDBs9sr34UaZx5RW7L5WcBTzhgz+LJmUEuwzp/leHWpc
X0bwfCOWJjT5FCHu1eOXiYDqpQW3NU4y31kFJZZL0gB/TDWhvKkVKCiSr6GV3KK2HOx13fucTW0Y
oILFAUk5BSnS/Mlfpqw50K4Fj47K9qEUsurlHs9q4pxHHsgV6OQcv4F3jpSqp4TySCw7vm1ygkW7
Hkk49ukZ0REACHecr6ac7pBmrE7aksU8ot9Czm/KpCMRNJEUdzfkspDGoXvnjsIWUehCvFOMXGBU
jJWGp9nwa+SsKY8N8pl3Q88uSbaerRRL41NgNX7qc4js1VU2CyUPJWq2X0cnPGgBHZjxjkLp5C5G
qgyLvzxpXucppzX5l6Il+g4rOVKO7uhdu1sUEUe1OPBoaWGUUjihwMX6kjI+F3r4PVzlSnfjjxUe
WU72idjjr7CDywI0IdN9r6aTA0A8BYXCcu1NipTbajQ7sSfu1UDzCqAYdvRBoEV6RPtxhXalLvHp
b1b+T3DFA8EiNqQF0S5dv5ubMj53jmjfOR9bIEH3+5CRehfkHDXFLopa5qd5o1HwcenM1/Toz9jG
4B4chz9+iodlJJiz0e7CbSFTN7x27lA9zpKhYqkB6c68Y9FrQdu+CLbKEbZNkrX/lxWaocuRyMnC
x/HjBYuRxW4IlFt45bWsVAEiXng4iAqGCqarMk29gUrrLPCO7gRNmuNsduvl+AIC55vT1Zng3tiU
W9QRoPdgyJrx7OPbntNclnEHOEJMuiu4nWzfLOefS+8S/DgjNSdVhZOcvshFHBZbA/QsiumM0lgJ
GB2dlyWBV+jPSmu6/79jlGCbuHrx4WwyufqchInBGgi9/fHa090+5Dv7NZobLO7kqKqDPXgmHJ26
ICZOFs0A1JvmlWW4oD5UQ1YP1cHr8Xl9cCnxrYVvO7qpZVzIJVhih8CBqsIz8PTJBpEg7h7tzfPM
pnwMVMnykYyELc3AalPCi66VpGBrDW+zT+7X61XHY+LBuIBXJyo0+RZNTZvo3sXhDhbrPga1UDcr
BgGT5GrqyszIHhdq/BI1fWmqMwhfuHEOtlb1goI/WZ0cRPDWebYCzgyjq0JKew2ZjVnPMOn8mqFC
Z4Y78s8SPR8L1BO7eMwOozV/gS+TY3BYfyXkcrkCSkeP7xIdLxUnmZHqdz4ci4bn1wm47w+AQmiE
YDVpYfKVfHwVQFXmYLbaszj+HOggYOxkMSLHNlSofiPG6ttpkH089XRD2X4J+YZ/IkntidrV9UGn
v0XD9rW01cfvD4cJihR5pWK82312VJFESgQTELg4zi+MSM9oHD4ceZvy8AUAzL3wHejKfK+EXgfK
bcHPOXu5yZYvYAmhACV4Oy7FHA3qh2Zx83ND8UPLceZ23vw9VCRbsOIrZOMzMSJc7yWCLdT93G9b
SdIYFd85rJbzFok77ANRc//9NFfBTOvSI0uTqjblVvCCrlyBvsn80m6WhZK/+1OFmQvArxMc5YFj
O7wJT0hC9JNUndwqD2coNsYuOOTknK+NunDjxgCXiEqpUKyxgvWvq14++J6XDILeX0vpOprSg+Cc
NL4O5hniWql8ETByqWgPS/k7mqzrbOnOk5WZC/BDmYABdib486xCItyFLN40Ejt6OfboyT9tlTXg
vT/lksgKhvYbbzGSKHYDtTYJvWb+1Znai/qcgoJNOenv8FP9ZcuqAcyAhwtE6EF7im1G0S9sQMgp
Lwo7aL5XWnp5WZgH7Bkwja/+tzhTFV9Q7Swb2JBc0yMz4k+pwZHxJNKIg6TM30OtmdSfu1KQkM4W
GNSa6mSABac+M8oxIdUg9FE/brsXVP4+QOASalmKoVF3qW/DZsZOZFvqlhK398aIGHY6DL6YUNfx
zZ7GdDySXHRduoDJcr7Nbb33kGez3teHXx4k0DjOIFOrMxVG6iRm00TMJnPLNEPyOu/2lFYvNUjH
YksKXxry8lpSqkCs/ld0aWGrR4uKkA8UzHuwyusNlV9h/LuuDzoozoe1hsKvEtbcMN1ZTuJQblvl
nKAtj+suWKWJy0Nu5R0MArFOk6rQ+Midjsn/sIgToMawGUhLWQ9Qsi1gQTDoGtThrEag+ypnvYEb
ugtBXsVMX7ehud9kde/EGCoLOFhqWSfKK2uObAcYmj6fAMTcf7NW6yPNpm/anC8ETDXafCHujQvC
EhYUlicXZ5zGYNJ+y3wRhRVCi0xt867tR7YBgbenqa8eVkHTHTBb28AlLfvsw+ivmTRfNbwclDuO
rP+Y6FYrqn6JBMzIIT1ZpmI9JQ/mRcZzCu5oT1J6e60y5d1xg4/w1f8lPdwlY+f1Ydk8SR3aTL9t
F+cqSgvJhozmcbLhr1R1qwirnpue0At1nFAeHENQO1lrDUmomTq+6v5oVxQe0nsJKzCfLT5N4aEb
MvMw32URXwkQ+icwj5IKxbf79dCw7zK5e7UtREAlW11Y5idSi9c9ZRmSK3XD+RQykBbAhlZ3KnyV
wBT0rnH+7d1wF4dvLXvpngaQOX8iSZ9nMOnlh0m1Dig1UN1Gd/al8+n6eHMXsL+qpGRNLB41Dq27
zOzc3pld75xnfCHDuBDIBG/XzRr7pClNoaD+GJzZdCPMyF6zLqKS30zQGWpx6GTKVbUVmTakLLir
X+dY31x0MjbViqxRbcoF2bTkL42jiGEw+ycycTg+gPparlE9DjpAtq4tC29HZWat4Pj9ZT87EelK
z/ETe3orfzaNd7l6RtOdO1hOpWHOyuqciE7OLitVRVuhUgSO0mWsPaMwzX79YnBGyAjKZ22ksNO+
yc/YLb8bBAyVlQgwZtOk/C619x2Es/dVM3mwwuAWfbu8aV7umRE/TIQtXPlUivbPWEW95EjfVFxN
s8Jg4unPYUNtHxYPLAZriYatzPtHrjSWcPdBlMvvuw8wwuq/V1k2/fV2+5E14a7RWAqTabDmtPKb
qxQfeUUhEiEhn5l59ALQuyu2HzWew4GjEMhrdYqEPNXWjcZCqpA+EhdglmNyKUzh/wAPsR//tLGA
gDq0EBesa/4CWEhtAY5CLZNR0m7NMrpGmZP8mDzuU1VkQTuaPVCCp1r2T8VxMLlN0eSoZM5ye8iC
6MmEV4SVD55SgrkvXX83eqWIUS46lSnELFdFWiYX6w7IKX304bC/pQJQZCfnzC8B+YRXTkC63MBb
g983GkqXw5biyD5Y7knop2tRNb3DlNmxrwkwB07o3wdpdz6n7TC1Ga4ii7pEPOc2S6WYx+jkR7Ty
/zH0Ol9cMId4mp6q1p61YOzLJgjGw7deca97pwJKYsrv8zeJ1dqoNSQp6CqXPCdwV01pxqwY3Qh7
t5cIoXAwPgto+fvc5A/Zsa6CqMkzKJ5aCTRLU/YIVjEgic+wuNwwgDw4re3UbGkefg3hT6IHtg/y
6ry0MKR67GMVcCh1rv0ME/5P6xV7NIbk6lxHOxmEs9MXQh9EKNsvzIm1yfdA8vXV93DY+peQEz6i
e4KO6Vauii90sG8sFZPPjMxe2+bdVnQQoZSH2kgneFGljfVFN9dAEyPpeyQ19697nNMbkIhEMpMa
FxBsBR3hHXE2tqYznAGFUVBpsAGbO6DyTZe4mVEDanjLzWA9lL3TvmTvmbExhy4HVRQ5nT+r75TP
tA6KsM5ZlZmchiN1INzz/Wmq8bjWUl+dIcNCLhhRSpCnh4gAzyFiT6fd5Gbw+N/2fSLW4XsecqVr
itxhuZgJ0P9mElFfSaBe2mdMZkyK8gQM/7987pRgJjaBjPX/mD0f9/DSKyz6FnToB838H8qOCXCU
eGByfBBig64tSc92PESOYGnftxNBRUonk4gn1Kk98pJzXWPqFwxltqAP5I0o7RyLNVVtSuzqKqYG
jjy3/eJMfKm36rT1kSPL8xOYqVJdbZovFL/Lwi1uIKvcJE7iG/zm9Q+N+yLAohghD7I5a+EK6ahM
AocPT1Jv0j6Q4s6fTbKAxMOpo8An/GwqwfFQN3qKLjRyLdR8AYvxKDZYZ4sgN8/XDxhn648ki4/b
TSDmSzoMDCF4LOvz/5Cu2reBXYJ+BkaeKjwcL7etkbreYXf/U5rXhI7t2o12W0JT8mqLAytNHK8g
rnQNgUmKfS0kRm0a22en88UKPK1iPjE4mhGk13pIR5ncxnCBFEKEChqGw98JmxGliuYk8hVcdiKz
8HO/vhIfI7I0cF2XnZRvVvmr7nY9J5WCIggWQUwxNanj6HcfKaats5/vQvY69lpqAViVTZQe/i3R
fVHaCSvMnD/KdeLjhao8zcKA6j3DwhX58IcZ1agCshfweW5ixvgYE9WKPr7ZZqUVgOW/iD6ZF4O0
6F9DEgfA1NxJaJ+kEDw7aon7LW6iJhfwc7ChMUwfbvi8QUWGYTcvZ73kkFnNHcMTMZjGWwbDrQ+I
BL+IRJONVZHGtrnIlRuusFe341Dj1cOVSca5lFJsLs7+ygoOCkjghKGvzJ2n9MAlwwaBEx9Ec2Z4
3h4/N+tVMDpKpvqvNjeeTDn+Kj39Kr7otDUMVYyTFVFEhPcvs4oeWQ8rfKTiYE2nz36Xa5z+CBK3
vRBtFtX92Y2jwTKs4Ka0b2K5LLE0s0Af+Rv5+AM5gKwd8vgIJdehyn91ltCk9QCmR5ztK8t8oTSd
EfrL6zjrctDxlxZmuhhiwrBofBVbxED5CFuiPxEwuy88LnOmLGhkIroalU9hrCL8priAyl3xNCLb
O177GHjGHQYiRqO3KJmQ+uBqLS9ZgUW73O/aMTZG6Netm8n4wAgsCmVPDIhXC0QEbeh8dQGiBTu3
yYewU9T3e3++I8QU4jFRx0DnRaQ5DmnMORg56I8S0l4B98cSeuQIycI1mEIADXHQz4POlhCW+CLS
mWOLfCOfKZ4z9T+BWI+Z14bkntqZXWyfNaUJFLzXX7cFL8lU/C43w2bqH0iWiPdFVNM3ZPVkKf0z
4LHV7zfqmjnrsi+LFZMyPky1qFOJtHf6D0r9ALsegBF1dJ0Nya50F8KPZoFFTA+bkdGsXzTWQ5T9
0rbBWJLSbJH2+OOGoAu2Tn1iS8jEOgasXC7afcFOZlqObf+T1m9pTHB40Ijj40bXusopKya6BnRl
9VcaVF+KqnAbwkELCnl5grQyYvAfb2C9/ci2q0c/N0CjfeRwajk7sIoiS4ihVtL14NybKNLMcvO1
f6lKgeUD7drreVE2iglQpnTHoUbTwkp1P7lXsJeSRwdcj5nCOjhddaLrCdDvg/uY5eJd6qCyovma
FKGNxLGtXo4LlStoXkj0mR+qpuPDRtnsvNCTnoTcPAjcHOKoAHmmvUvqxdDGmEEOUCKOhzAcDXGV
YU6/TpEZlBdfnwb6wUgYxsS1wnJhLhMQ9cIuEdjYTgwkRlMjh5JeJBO13oP4bmkolb0LP4AumVGh
JK/d+uulj0Oo5oh01GvQHONi4UQ8oCBt92MjRDJodmw9JvB0U/2pme44MTKaZLzw3DvmNztjoLvx
yZ2kcjExNAXu+tZbLvEL8VUxGS3k4YBKkPIhzZ3g4vwuwwOGyMa0hRAZDhI5JplMnKtcqFZ1YWoP
uLpxBUqf5X86IL7QVduxc8pEkoV/NoZ+uMh2XnTW5WKMRqMGbzuExWVKZ7l0jk9xSB10j9cYl2oV
SsVwGfUCPuKx4kzo/Fd25qDI6C5ConKf0u8ZZBd3h3sLhyeSu6HHedfW0ngACmn1ZBrk04sOxmm0
PImdWJaaBT92vuZtRy6yqGieK3aA1aTqWwCSqqxGAxSCpjsaLFEH6ZEKxisCCFYusHTW/vWRASUG
j7po3gGFCLlSbFWMdBPIh23qtn0yMBei3TBu1SbFOtHvNygxuO8UtEhuBNZGdF//N+bDoRjVAvde
LWqAlec/oJroZwXm0ixHvU3Ss0RMIGT9jTYDRfLmR7Ki6dOlH2doSdWjVtn3ry+QIXjysujAg8+G
uJSNkoOsmTMdl1x68kSTe7UnPJXU5UIgKqPy8W5Q9DdwElUAp8lXO9MRiJLMstzzUtDYDKJ3qMSC
p9+8BLEgBuDnDlSlys8l9LXMZawCqH6zalT0g720zjGxm4Ofam7e2CHto36HCeBPwU2KJFiuALND
f7ezJF5+YTCVtMNV8n6DxPkfsz/PvJP5MwABwwThqXE3MriOk0s43ue6FU5EcfL0vmhkLaRGYwvV
fRdIWFSq067OxMfa6RiYAybAVoAAcslc0pf1oUTUFT4DS7pXzO4rTwZr7GxIqVZHIKGDlIvRrMQ6
52P/Ntgi1GXb26MTUWG7j4cgDDj/BEPph3wU6lUzi80v/aTrniNkkAK1ylZUoOnJBDtfXXfaG81K
MpM3gXGsRLK8//V+hczdz5+XserDEEKzijwtX23z+TVpKO4b7jFiEVn0EaXoCx3CAKNbWI9hJm65
wugrvMGHed/vv7b7xKTy4VSdBc6mffwnUp4gt7D3RLNtMp+ZfO5irlSrj0Ka8UHCCQAB8SlvRK3g
nMnz2Hca3OvIYNo1yowhVtjYilNVRvAr/TbnOVeSUKYs2AwUQ9tsuH5Uge8EsyJUApJWcFExnInL
zUoauqMOmerYahJfOnSprmZbprVWaK44V/CbBGT1XNEYhkyudCcu200Ca8SjIlX7gE4PBnTJNLBy
MeQalHEccnQ9mVgqmvtjvlHlnXfHC5+ItdLdY2JKJCyxYaElUDhxz+9emLCGUpYmY3yC8kg10zSD
LVFpDMzh3bJXMQ44TQhCyZcwAjSSxw7Ujrn6ddvbPF9NJeJXo6QNjvB3yfS04DzfLVXXSUG/eJv/
eAebABbd+hip5kYb68oUlTmess+2A1zd2+Yo2cstT9EoklOF5DEjiuBPJUgYFR480neWiy43aG1i
dlv8WM1Gp8oLhVl/CmVeuSYgTZLR92/UWDfTtJbz+hPnzdqbs4pT+t59WAcjLjAf6+A7YspESrev
9a+57REB6Okzj7ZmIgobs5KYRXxOUz+7sqnjVV0W6OI5Agv7PP9SxTlnXVK+gkQ3U1Bw+Yj2tlxy
gSWR7aTqksMhYUnFthxec3OmI9qnfVMZ1HxTOX9Ol+HYhTog/RMIFmDefZR0i13UktQtz7vpztXD
CKsZaVKPgqs6FCs5Td4TqO11c4e8nqmL67jbzGMVTKrIStYyRUwoOkrCpWUuK4yb23zOPSMSUXE8
yTdj8mpMkVw+aDse477ewSk4oc/cVnxWACT5vyLm9Qv4InOKYlewG4OZBrcPDREtApa4Vs8We0x+
KX4dJcfuKvO+4/Xx0pwHJ5OH1UYhrP8w8fb1aLUjm1yzKWjPCNbf5yKDlXkSSntX4567qfEhXmn5
DZbFOFh/tXYJvq8lNq4wkhshpE1gYua03QkVe2jJRnxZf/aeiIYVDJvSMf6CgB93adbjDcu8kx1p
7/j4qdbdivlbiIxS/6KXMlYTAboQzxZRuueRKIvwhYwHVNfv3Irj2vfgkh25k0oUC7/fwg5DUkz1
amQRdWejgCKqRZ6IX7iZ820J0vqiK7MJhqD2YKhW1X4roI/CWNA9EFL9pO0HkWcQ+gb9EpFcccE6
WDoNDPtcKpUU/n1MGP7Jq81IvcQlGrkzIqaTg3Ly8pDIksLFc4souhP3ebT61UxfQa91gWrJ0BzR
X4dVF5TtSbxrxrxbNxoD9uzMRzSwIpMeEgO2Yr3J5BJvxG5Z3WTd1VwfSEX2Y5itfl38dGe8gewB
w/xtvDn+STtvTJJZ1Z/S9gqD0EnGOMmZUhiFUD+BNLGfIyWGrYEzhCaAQzVNxiVHVruj8o2NZZRm
i+hA/GzMtK9Bo6PA6Nqe/MJmdDQwwvS+Vjn1vmtA1j3/4baBAwA8TwqIBABHFIYyUcHwGtM47g80
nfIKuoJUJC+DMFh4qOCWtNZb5RPZ/L6v8jChI4gmpqAfTj1nM9HS1wXag5WPbB93j7zXgwJGHV/v
H7l5ENlZkh/aWKHb5xC3sHOL0UIjYmKY2Ebxi6R0Qe+HxTxgqxH0MLNCo3ObMHZtIFlEjSAm4Kvb
KMZDxq4QuLt0sPuecR/L/uPxcwchTJBbatXrqGwwXt/Ud2B70M2QCankNSzpie+uCNDPtvlzss2H
mBnE1n42Yr7viNaHPCtZKgsfR7abSf/oDDR3iq4/d+2ppsLV+L63d0V9sMYnL9jKax8ppgUqIzuR
Sjg+DfvNdyNAhbK+SQsotmbcdz64Vykv08ejx2yYgrDPHWh29T/g+V04+lp2Rh/uI+MQkgfJcUr7
O+9J9DEYlKyFSAvMZmg0zMpN2vxqkL3qNMv97yVjWL7oMx5KnjsX726KZUZFV3jJq2JmoY9K3rHK
pL4dJgKuGR66BjO3kPHcLHWG3WYjotpu5pSS2c0fJAYfPUorvxSe22ElekFfh0HWJShhUjvY6zrY
zKw74j71rf9t14z7q8Kpimt8kNTkBKdD2VsQ3vdI/ECkfTYnt438aaiy5DV/Wj4qV8lAp48y0D8x
+AuNsnTU+kqNZ6Kco8glRejQQUGjgFm2V/VQo7c6U0O/qrEJL2q0boQcWIkXUKCInHPTrIAyqHkR
CzxIegVseuZEWmc3yLgeQzdjIWdhaBGnHO4TMjbT/LrVSgYcTsCnriULEJYcOShMnObDtzVjriwZ
m0xf0rs45PIZdQ1RhMmivgJA+Byt1883Q8wauMYgR33InbkbKwGC4bAsyJurE3i77hEb28gTNFTB
aWezEgAeHhPso7OV/Ju258dJvQp1OmlecTqd5P9a9BuB+8/Y1HNafGlU9wRnDZYwf7EBPh06OB/R
hwZCTyGUVhWrayv7gCGv4A/tPqRh09w5FcA6FPVpj0r5USeq/HFJVnk4If1AEBIOevg9W+FlNF+C
lKf6Zn+G30Ab0/lcMMV7d/5b9vGHI9dFxjHNCOrLU3QgfWxFzywYvmQfLdU1lakoukvO0VZ3YTVy
0Mt43ucDO7iByuLkJVXToE/ONgZUZqEJc8icxR9DV0XaZLmC15oRQD6mStlSeJXqMuRZKW1EAWB9
NG1fI4M1TJ/aoisbADlIdtEhQ9dpLBYkIsBUnqaV3/wO/L0WWbxzahZwNoSu7SKVF+Kanp0/vnoq
veU8jvJ+5+k94W9OmUgIlu3bDeQd9S2Op6ao+QrWPrnFLkiaJWRZBiBizw8Eo0X9vOcXzTWnh/XD
QKFMkq4h+4ZXfyrloTQHtH8CezlAmHFmV5MNkMpGDgqCwMaht6/ZRjbWTv3UNPwwx0BwK0j2V4/t
i4BNDtUR1oN18gMau5nd4wXeJnKgmfyoVykmy9VJtypH1t2GvsXRTbEcA2/+BvdHnkvPCzV1O7Mp
HXX3hpQzDVU1EvNZDb9SF1zHEf+iDemqYjCZfC8zk/yapxturGBNA4xUjwMALGmwSwjShgnZRfqv
AcNVMmcn+RJuh/w9U5qOwZzWvw51Fpf2N5evEM8qIhZnDCdFYTTWpYm6679wMskaYSBdel/jjZb8
xLPYFrXjcx4hkmCaRpB6lDoqtLsKAjyX11UNQaT79vg6DXy+M5rRjWahY7a4wjSpBun1k5EkOhq+
zM9zE7mNh4qHkPDvEcb+nGJKoaPgQ7K3VI4p3D2rod8z5yToIKMgvKMgaHZ+tcXGYYr03HRyjpcK
A1R90hmhCrc2qUNZXsHRqjsfoERvpKkggtxuQhtgmI2CtnI+bn2sui2gypNy5zy+reQEn9MM2ew3
P2pdfI9vGya4oU+q4Rb55k1y+DoNBR5rJ+6Mm2C3aXSBZm5JafiE9K4kI3wpgxYzQ1HFSFqzgruX
o3/PT3zPXKJe4pmpLNoUEhw4q+yeu4evFncLNiggpexlKFn+nbx8P8Sf0GW3vNUp6sz64Yi+ebDn
c3LGjPvhT6fQbkPeYnkSYvTq6YLXVvxYiymh/0q/IkSgigVjkUmx153w+wKAdmA72DLDEyniCLAu
bcvehZtFxF+YzlyJ37Py+a+I3ILQ7z7/+9pJiF1G4yTiKz199QKKvBuM6YfdP4jaYSOpEbshTbpk
wXJ7xbQtnqX83Ww3z2H3Kbi8AX4VjI706ziX8vbTYq5juP0dgaeMElO5Mj+udT1frScqgxNV9dkJ
clWklKxPPjJI/x02VHiNJ1iUFL3GL46upZRzpFe+7H/ZgWTiYx85md1MKFIOSX5mNn3WX370LJp6
mN55Lsk9TM3CWpQMCXOsbu+sO35rc2rSbtPcQx0IsOnQK9YvlknBowrB36tcIQYuJLFfkGPOjPKT
E+SkbcRbTTJHdaYNDgnkxtXcivzfE3I4mc7e6goRjY/tRNo5giM+Zvf+vBhN3VAyVXprWcxVnIbl
GdxAU1at7I0NhIf0E4ridUrhgNja0b+m81A0uAdexRFBIPbvfyvUbo6ZOtCN8M8l3v77OWuLhaKy
zKZCWL3Aj2XzuDVEzcYfb6/R4A6TMGSvMlLcAVrgsXwGFpdHaST9Y+embJyzY5Vv++TdOhcgHuxm
+9ezWYhZGdHA+vG8A+ExFOECK76IAWthDFVo2Bt6xvA344fT6cw+vujyeIbyTSvWuGUrdTHPtkHF
CE9e6mgl+EmP9La/hnIYA52NvcqxhNFE3QfhHG6ofeGJWdhdonY6fs2bsjtDip9J4eIJZu0YofXT
rTEr7OQ2GKKzen/pbKpT+g0XtbOAzpD7rgw7rw/0X14+NsTfiFkti4I6j7SQJsJ/0Jn4BT5O67F9
B/r568lOapclUQBkENg2yztw9qxdUz2QXUKOKQFb1ANgt7UWItkoB8KMm52kMeqYFlubAH+WaOu6
IfvL+4KZlVpXdQEmRaa2XVu2oKKTj6m+L1L6g8Tbtl75dOySVig8DpQSGv9ipJPE400mOo0D7i1V
85m/KRPYmi+91RsfLZKPDtlNyvRA7OaouDzWanuNTmTS8737NKdDs1vZtpLtckhjNoNQs5fBosTf
dQ4nRrckELsWDn7pVoK1esfzzHBdC3f1tWS4cUoMCFNSHAGKRTAS1cgDOPcZnoQWqF7aw3I6XJaQ
Iv5nj4Rn89ITUBmASb4KAGEWIRAL+1zSCR5DKK91IndV1LjGe6FHE07BrRWuz2mNSOIiQRHz6FGu
j2JhCaDry5b3Qb6okD6kcVJfK7MjeuIr8au2qwcf1kzVQ4oQ1HyAHomZGuM9imyS1ytar9CsKwQu
bEquOYYDxByRN7L6d7YoeX+/dw3vcyiWESzPFiCVPVWYC7Kg/vuPEeqwzpjAg62Xp5TyEx8w+Ukw
Mem2Vb42yCiC9OsSj/uoucyjAZAVxSaBbU6+fBDBTBTzIjyxSC2G6PRH8HOUUwYoREUC8Cvu+rxF
niR5zFM3qrcTBbV1US2IH0VbgtaDotaKI86txsRGcf+XIGnc8jBXIMGhPiE38b3TNItWs6UiF68m
E+cNvC+1KH2ocsolAFiW4AJPo08a4lD2K1alNCKeeo2YIiCL31jra5RptvKDywcbjlv4OGs91uAn
EM+FYxnOGMVg9pPoDD18m+QX/d06mPs8h0Ew6Y7PG+3LlrqWoEDwvHvxRZFTKZ1SH7cCINmapQT+
QaBXL4n6+8Wsc2+ZaqDz8LI7f+laLeMtRwKDuG7yItxMex70znqFhfXpUpNgNVemKjqV89aqOAjP
E8RokGNvOPQ8g5pO7fiU2bQN1cQKWk5JIj2u61M768DB9F+7FENpGjoBNMeDbeJ/kv4xBpvlCEtt
zi0DRkxURlnTAc6NZyPTlgsj+Jg8IwcvphLtYih/QVXuL1n94aWmJzADUrYSM5jkWJT3sOFse2LA
OiMvdggXpVhcsh5eCaOVdveyubnOJpcVVGc6uRU/myi299tIWdjx5A/coaP2Cqhvbf9FvKYPn5Vo
inznfADAhpQb2j4ZScR6fncn2CXVfsxxYq+nZnXwWAeMAkVLoCIHjCBzn6viIBqnntbPHMRTT8AF
rvNZ0LbL+OXLrVE7mAfO/+OMXIg+cfYyntuQ6eVXOBAmQ861RfSVvXrAUk/1IXx46wEY5lpj9WMU
Le5kN2Du2l14N4YUmOxskXPuOWxkx953J2svbvpYzfnkc+I5z1EMpntTiditMKUsoBhtizvV10Uw
D20R3m+a+1y3SIeHH3SDm+9GtyBj3jVU8733KxGru80EPLSavl2rhAFJQSJw2EymlXDzQjmVu5cD
nyxLWKiD/MjaMzPawOD3v5W7GE/IulFEwB4JW8CdqBjlyx9Kii2rsje72IsZaN0lSvGJFsrC5SuZ
73mESq7TpktIb8/G7A76hhn8wk0jiu3nGh0cULOPyqGeHvyoXIshdHH//Zx72LPuw53IbwDRIJcj
f4gTne7xKKJK/qlq+/mqm3q2SFlUODMDBKq7MjWoDsFOqDnlsTutSIi0tBb/5NtipSPnjof9ypac
tr5j8SyPyG19E9MP6HtmtuRthChDpfEayWjWGBhvnrwgqqpJNgUhjDgvIjw/I2q4EclGm0ITvnPz
ZGRY7hk4En5c1xbhtyqfEkn2imtRml31tl8FI4mybKNdY6EjhACjmAPgRGQrPdEHoDhQNJbHhxim
WWigbTSc6FfUpqXyr9BG0gZyyxx2Iq0Bj+XRoDemCOofqFk9+i9mlbSWRWGfl3BWYR1Z/fNMxSim
p1yqggdFNcYJhXeG4o7W2ejy9u67wTQxV4PZw0ZsVPwWXu986Wb/o8JE0HXeeSERA30Cs/bh66ci
rwELFlfvh9+Lyla/jxtTqlxinqsPq6iyICPtUWguUwTMthPfe0Sgb6inMnrMDVhYlyfsIdwWglcj
tt26jnL2ITeFGzAtoo9CsX++KaWpun0OpRByWopi9VQCyMxotVBpDQCaqE85c9lZT1Ea1vUNq/7i
e9aYuGgZRVL59Z/v1q2pg0H/4olcC5QhpcpQroDNM+GRhQ9ObX31j9+xKPIOGwPgGnwHTFPraebs
rxiuHdf7V33SKMKqx0G7LkUW4MBBfBElZRMXEd1UMGUfQqE4tJ6mUhH8qXeWvkO3HUoAUn+wzuHK
abM3wVteKq2xvBxvTZt6BdCNJ7rNQKVFSDanurwW8ZMnRUMGLZC4gPW0O5peZ8iorYA8Ku+eM51p
glDV6gZLu+0TzX+x5wkxCZaU5wvjSt6Gv+EOG/d1rEB8KRrDkHP2fRPAilHhKQfC7/aLWdAeUitZ
AXi/wdFJk4922fAksQvK3DmirKV83b3wQIMfH0YjJKvMNoktFWv9N5zLAuCse1O2PJbIZU5iFZHV
ZLBOgch/AMZ2NZDyGYCYlLtBgL/NjF9jSLtnukrxa6NYUB//YgM6QrucG9hhqeGJLxbnyCBI/EzF
JuOuxAtGy4uSJlNMR5lhx7E+AClhQWKorY2pM0ff4OnP33pWQj/SKv/zppwx7QCa156+2QyeN2su
y39WwX7fkenCm63JOuyFyFlJg/zSEr19JWxb2ygzMBJDLmefpt/gh6/s+YzmAnjxsXuF6MGlwoVT
kB7Ea/b1Jlod3PsdV9PXK2T6WNfNlv8kv09DSn29WXXHosCnMYbilZH0WFfPFSIGcQLvRI/W9hoV
HnyYUpNsz7jreM+ueXE9PYekFf/Xfa9F0kzbNWMFvsmmrofYXOV4inLllraeJl8BX1VWiHDNimzL
hQnOzBEghZ/f8IsoLnasyXVpFXbcFq1Xs2F2shAZHZ1wGvNEvwYWgHmo38zzsR/TAKmTYXtdj8N0
VLGa+RWzMIWpro2TkhMhrwFV7koyPzCje2Bt+yzYpp8Z/lIE+4N3UU3kM1+uKaFQoRtCSjvvbBT6
lEFI9NcuCLo5vkNxkOLhKd/uwQRJrJOiKJ85ULq5mtPVuOHj7lBtgQUXyFef1Utzao/7VtZr61Ty
iPzTDWtfwYudxWodZ87cizj8A7m+GTH1O5voYMhxWXihKJwT9SaOMdT71ieiJoGrNREwHI3oB9dM
lI8LWpfslSy5eYHrJ5DFCZJahIwgzxKaUYbiJfywzppsKugOynxjyc6v/M6I1NVEVDNgvckmdFFe
cJopni26Ym1dNgVbtr1OyFQQQZMwi5MC6/k4nHmpQ+R/NCMvXGCEs/4kKqJJVBw2Kl7xYfhn/MwZ
gTQ2EJ36WuUfZhslbGjUB/uEZxhHwVeSfhf5q6Ev6R+0XsEYvYzZO6ZQ0QLzOqvGNkkitKq3JdfF
pKa6gIwD5dR8/hfLcmDtGuU96FS2dcz24WmzcDJNjbgZydFu9zkBfiD5gEX/KQ3HsAIWVc7CduzE
pgmRZtUx2M81
`protect end_protected
